
module part2_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   N46, N47, N55, enable_f, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n107, n108, n111, n113, n114, n115, n117,
         n119, n121, n122, n123, n124, n125, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844;
  wire   [9:0] a_in;
  wire   [9:0] b_in;
  assign f[19] = N55;

  DFF_X1 valid_out_reg ( .D(n844), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[19]  ( .D(n81), .CK(clk), .Q(N55), .QN(n821) );
  DFF_X1 \a_in_reg[8]  ( .D(n119), .CK(clk), .Q(a_in[8]), .QN(n805) );
  DFF_X1 \a_in_reg[4]  ( .D(n115), .CK(clk), .Q(a_in[4]) );
  DFF_X1 \a_in_reg[2]  ( .D(n113), .CK(clk), .Q(a_in[2]), .QN(n803) );
  DFF_X1 \b_in_reg[6]  ( .D(n107), .CK(clk), .Q(b_in[6]), .QN(n811) );
  DFF_X1 \b_in_reg[4]  ( .D(n105), .CK(clk), .Q(b_in[4]), .QN(n808) );
  DFF_X1 \b_in_reg[2]  ( .D(n103), .CK(clk), .Q(b_in[2]), .QN(n148) );
  DFF_X1 \b_in_reg[0]  ( .D(n101), .CK(clk), .Q(b_in[0]), .QN(n843) );
  DFF_X1 \b_in_reg[7]  ( .D(n108), .CK(clk), .Q(b_in[7]), .QN(n842) );
  DFF_X1 \b_in_reg[3]  ( .D(n104), .CK(clk), .Q(b_in[3]), .QN(n809) );
  DFF_X2 \f_reg[1]  ( .D(n99), .CK(clk), .Q(f[1]), .QN(n831) );
  DFF_X2 \f_reg[5]  ( .D(n95), .CK(clk), .Q(f[5]), .QN(n825) );
  DFF_X2 \f_reg[9]  ( .D(n91), .CK(clk), .Q(f[9]), .QN(n826) );
  DFF_X2 \f_reg[13]  ( .D(n87), .CK(clk), .Q(f[13]), .QN(n818) );
  DFF_X2 \f_reg[14]  ( .D(n86), .CK(clk), .Q(f[14]), .QN(n827) );
  DFF_X2 \f_reg[16]  ( .D(n84), .CK(clk), .Q(f[16]), .QN(n829) );
  DFF_X2 \f_reg[18]  ( .D(n82), .CK(clk), .Q(f[18]), .QN(n832) );
  DFF_X1 \b_in_reg[1]  ( .D(n102), .CK(clk), .Q(b_in[1]), .QN(n807) );
  DFF_X1 \b_in_reg[8]  ( .D(n841), .CK(clk), .Q(n812), .QN(b_in[8]) );
  DFF_X1 \b_in_reg[9]  ( .D(n840), .CK(clk), .Q(n813), .QN(N47) );
  DFF_X1 \b_in_reg[5]  ( .D(n835), .CK(clk), .Q(n810), .QN(b_in[5]) );
  DFF_X1 \a_in_reg[3]  ( .D(n114), .CK(clk), .Q(a_in[3]), .QN(n804) );
  DFF_X1 enable_f_reg ( .D(n80), .CK(clk), .Q(enable_f), .QN(n814) );
  DFF_X1 \a_in_reg[5]  ( .D(n838), .CK(clk), .Q(n806), .QN(a_in[5]) );
  DFF_X1 \a_in_reg[7]  ( .D(n837), .CK(clk), .QN(a_in[7]) );
  DFF_X1 \a_in_reg[1]  ( .D(n839), .CK(clk), .QN(a_in[1]) );
  SDFFRS_X2 \a_in_reg[9]  ( .D(n836), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(1'b1), .SN(1'b1), .Q(n121), .QN(N46) );
  DFF_X1 \a_in_reg[0]  ( .D(n111), .CK(clk), .Q(a_in[0]) );
  DFF_X1 \a_in_reg[6]  ( .D(n117), .CK(clk), .Q(a_in[6]) );
  DFF_X1 \f_reg[2]  ( .D(n98), .CK(clk), .Q(f[2]), .QN(n828) );
  DFF_X1 \f_reg[3]  ( .D(n97), .CK(clk), .Q(f[3]), .QN(n824) );
  DFF_X1 \f_reg[4]  ( .D(n96), .CK(clk), .Q(f[4]), .QN(n834) );
  DFF_X1 \f_reg[6]  ( .D(n94), .CK(clk), .Q(f[6]), .QN(n833) );
  DFF_X1 \f_reg[7]  ( .D(n93), .CK(clk), .Q(f[7]), .QN(n822) );
  DFF_X1 \f_reg[10]  ( .D(n90), .CK(clk), .Q(f[10]), .QN(n823) );
  DFF_X1 \f_reg[11]  ( .D(n89), .CK(clk), .Q(f[11]), .QN(n816) );
  DFF_X1 \f_reg[12]  ( .D(n88), .CK(clk), .Q(f[12]), .QN(n817) );
  DFF_X1 \f_reg[17]  ( .D(n83), .CK(clk), .Q(f[17]), .QN(n820) );
  DFF_X1 \f_reg[0]  ( .D(n100), .CK(clk), .Q(f[0]), .QN(n815) );
  DFF_X1 \f_reg[8]  ( .D(n92), .CK(clk), .Q(f[8]), .QN(n830) );
  DFF_X1 \f_reg[15]  ( .D(n85), .CK(clk), .Q(f[15]), .QN(n819) );
  XNOR2_X1 U124 ( .A(n810), .B(n811), .ZN(n293) );
  BUF_X1 U125 ( .A(b_in[5]), .Z(n787) );
  NOR2_X1 U126 ( .A1(n456), .A2(n455), .ZN(n122) );
  INV_X1 U127 ( .A(b_in[3]), .ZN(n123) );
  INV_X1 U128 ( .A(n123), .ZN(n124) );
  INV_X2 U129 ( .A(n123), .ZN(n125) );
  OR2_X1 U130 ( .A1(n512), .A2(n511), .ZN(n535) );
  OR2_X1 U131 ( .A1(n264), .A2(n263), .ZN(n602) );
  NOR2_X1 U132 ( .A1(a_in[0]), .A2(n813), .ZN(n305) );
  NAND2_X1 U133 ( .A1(n308), .A2(n307), .ZN(n386) );
  NAND2_X1 U134 ( .A1(n481), .A2(n480), .ZN(n485) );
  OR2_X1 U135 ( .A1(n483), .A2(n482), .ZN(n480) );
  NAND2_X1 U136 ( .A1(n483), .A2(n482), .ZN(n484) );
  OAI21_X1 U137 ( .B1(n277), .B2(n276), .A(n275), .ZN(n320) );
  INV_X1 U138 ( .A(n272), .ZN(n277) );
  NAND2_X1 U139 ( .A1(n242), .A2(n241), .ZN(n263) );
  NAND2_X1 U140 ( .A1(n238), .A2(n237), .ZN(n242) );
  NAND2_X1 U141 ( .A1(n221), .A2(n220), .ZN(n222) );
  NAND2_X1 U142 ( .A1(n219), .A2(n218), .ZN(n220) );
  NAND2_X1 U143 ( .A1(n215), .A2(n214), .ZN(n216) );
  XNOR2_X1 U144 ( .A(n219), .B(n218), .ZN(n194) );
  OR2_X1 U145 ( .A1(n549), .A2(n548), .ZN(n661) );
  OR2_X1 U146 ( .A1(n223), .A2(n222), .ZN(n606) );
  OR2_X1 U147 ( .A1(n189), .A2(n188), .ZN(n621) );
  NAND2_X1 U148 ( .A1(n389), .A2(n388), .ZN(n441) );
  XNOR2_X1 U149 ( .A(n171), .B(n148), .ZN(n334) );
  CLKBUF_X1 U150 ( .A(n360), .Z(n363) );
  NAND2_X1 U151 ( .A1(n445), .A2(n444), .ZN(n446) );
  XNOR2_X1 U152 ( .A(n258), .B(n272), .ZN(n284) );
  INV_X1 U153 ( .A(n219), .ZN(n215) );
  INV_X1 U154 ( .A(n218), .ZN(n214) );
  NAND2_X1 U155 ( .A1(n507), .A2(n506), .ZN(n523) );
  NAND2_X1 U156 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U157 ( .A1(n503), .A2(n150), .ZN(n507) );
  NAND2_X1 U158 ( .A1(n479), .A2(n478), .ZN(n496) );
  XNOR2_X1 U159 ( .A(n503), .B(n495), .ZN(n508) );
  NAND2_X1 U160 ( .A1(n485), .A2(n484), .ZN(n510) );
  XNOR2_X1 U161 ( .A(n505), .B(n504), .ZN(n495) );
  AND2_X1 U162 ( .A1(n497), .A2(n496), .ZN(n143) );
  XNOR2_X1 U163 ( .A(n434), .B(n481), .ZN(n475) );
  XNOR2_X1 U164 ( .A(n483), .B(n482), .ZN(n434) );
  CLKBUF_X1 U165 ( .A(n553), .Z(n588) );
  XNOR2_X1 U166 ( .A(n318), .B(n282), .ZN(n324) );
  NAND2_X1 U167 ( .A1(n288), .A2(n287), .ZN(n323) );
  NAND2_X1 U168 ( .A1(n286), .A2(n285), .ZN(n287) );
  NAND2_X1 U169 ( .A1(n284), .A2(n283), .ZN(n288) );
  OR2_X1 U170 ( .A1(n285), .A2(n286), .ZN(n283) );
  NAND2_X1 U171 ( .A1(n322), .A2(n321), .ZN(n325) );
  NAND2_X1 U172 ( .A1(n318), .A2(n317), .ZN(n322) );
  INV_X1 U173 ( .A(n143), .ZN(n567) );
  NAND2_X1 U174 ( .A1(n408), .A2(n407), .ZN(n409) );
  INV_X1 U175 ( .A(n572), .ZN(n557) );
  CLKBUF_X1 U176 ( .A(n556), .Z(n569) );
  CLKBUF_X1 U177 ( .A(n641), .Z(n642) );
  INV_X1 U178 ( .A(n661), .ZN(n666) );
  CLKBUF_X1 U179 ( .A(n719), .Z(n720) );
  INV_X1 U180 ( .A(n709), .ZN(n710) );
  CLKBUF_X1 U181 ( .A(n602), .Z(n139) );
  CLKBUF_X1 U182 ( .A(n608), .Z(n137) );
  CLKBUF_X1 U183 ( .A(n613), .Z(n138) );
  NAND2_X1 U184 ( .A1(n622), .A2(n621), .ZN(n623) );
  CLKBUF_X1 U185 ( .A(b_in[2]), .Z(n778) );
  XNOR2_X1 U186 ( .A(n435), .B(n475), .ZN(n127) );
  NAND2_X1 U187 ( .A1(n274), .A2(n273), .ZN(n275) );
  NOR2_X1 U188 ( .A1(n274), .A2(n273), .ZN(n276) );
  AND2_X1 U189 ( .A1(n180), .A2(f[1]), .ZN(n186) );
  INV_X1 U190 ( .A(n453), .ZN(n128) );
  INV_X1 U191 ( .A(n128), .ZN(n129) );
  NAND2_X1 U192 ( .A1(n217), .A2(n216), .ZN(n221) );
  XNOR2_X1 U193 ( .A(n130), .B(n450), .ZN(n455) );
  XNOR2_X1 U194 ( .A(n449), .B(n448), .ZN(n130) );
  BUF_X2 U195 ( .A(a_in[0]), .Z(n131) );
  OR2_X2 U196 ( .A1(b_in[0]), .A2(n807), .ZN(n365) );
  INV_X1 U197 ( .A(n181), .ZN(n132) );
  INV_X1 U198 ( .A(n620), .ZN(n622) );
  NAND2_X1 U199 ( .A1(n387), .A2(n386), .ZN(n388) );
  OAI21_X1 U200 ( .B1(n387), .B2(n386), .A(n385), .ZN(n389) );
  AND2_X1 U201 ( .A1(n189), .A2(n188), .ZN(n620) );
  NAND2_X1 U202 ( .A1(n240), .A2(n239), .ZN(n241) );
  OR2_X1 U203 ( .A1(n240), .A2(n239), .ZN(n238) );
  AND2_X2 U204 ( .A1(n136), .A2(n844), .ZN(n133) );
  NOR2_X1 U205 ( .A1(n436), .A2(n571), .ZN(n134) );
  BUF_X1 U206 ( .A(b_in[5]), .Z(n135) );
  XNOR2_X1 U207 ( .A(n435), .B(n475), .ZN(n561) );
  NAND2_X1 U208 ( .A1(n684), .A2(n683), .ZN(n136) );
  AND2_X1 U209 ( .A1(n844), .A2(n704), .ZN(n140) );
  NAND2_X1 U210 ( .A1(n705), .A2(n704), .ZN(n141) );
  AND2_X2 U211 ( .A1(n136), .A2(n844), .ZN(n145) );
  OR2_X1 U212 ( .A1(n795), .A2(n821), .ZN(n142) );
  NAND2_X1 U213 ( .A1(n794), .A2(n142), .ZN(n81) );
  AND2_X1 U214 ( .A1(n768), .A2(n149), .ZN(n721) );
  NAND2_X2 U215 ( .A1(n140), .A2(n705), .ZN(n768) );
  AND2_X1 U216 ( .A1(n788), .A2(n844), .ZN(n144) );
  AND2_X2 U217 ( .A1(n136), .A2(n844), .ZN(n767) );
  BUF_X2 U218 ( .A(n201), .Z(n421) );
  XNOR2_X1 U219 ( .A(n821), .B(n669), .ZN(n146) );
  AND2_X1 U220 ( .A1(n654), .A2(n653), .ZN(n147) );
  OR2_X1 U221 ( .A1(n795), .A2(n819), .ZN(n149) );
  OR2_X1 U222 ( .A1(n505), .A2(n504), .ZN(n150) );
  AND2_X1 U223 ( .A1(n586), .A2(n585), .ZN(n151) );
  AND2_X1 U224 ( .A1(n650), .A2(n467), .ZN(n152) );
  OR2_X1 U225 ( .A1(n795), .A2(n820), .ZN(n153) );
  OR2_X1 U226 ( .A1(n795), .A2(n829), .ZN(n154) );
  OR2_X1 U227 ( .A1(n795), .A2(n832), .ZN(n155) );
  OR2_X1 U228 ( .A1(n795), .A2(n818), .ZN(n156) );
  OR2_X1 U229 ( .A1(n795), .A2(n817), .ZN(n157) );
  OR2_X1 U230 ( .A1(n795), .A2(n816), .ZN(n158) );
  OR2_X1 U231 ( .A1(n795), .A2(n825), .ZN(n159) );
  OR2_X1 U232 ( .A1(n795), .A2(n823), .ZN(n160) );
  OR2_X1 U233 ( .A1(n795), .A2(n826), .ZN(n161) );
  OR2_X1 U234 ( .A1(n795), .A2(n822), .ZN(n162) );
  OR2_X1 U235 ( .A1(n795), .A2(n833), .ZN(n163) );
  OR2_X1 U236 ( .A1(n795), .A2(n834), .ZN(n164) );
  OR2_X1 U237 ( .A1(n795), .A2(n824), .ZN(n165) );
  OR2_X1 U238 ( .A1(n795), .A2(n828), .ZN(n166) );
  OR2_X1 U239 ( .A1(n795), .A2(n831), .ZN(n167) );
  OR2_X1 U240 ( .A1(n562), .A2(n127), .ZN(n168) );
  AND2_X1 U241 ( .A1(n558), .A2(n572), .ZN(n169) );
  INV_X1 U244 ( .A(n803), .ZN(n170) );
  XNOR2_X1 U245 ( .A(b_in[1]), .B(n170), .ZN(n176) );
  XOR2_X1 U246 ( .A(b_in[1]), .B(n804), .Z(n190) );
  OAI22_X1 U247 ( .A1(n365), .A2(n176), .B1(n190), .B2(n843), .ZN(n193) );
  XNOR2_X1 U248 ( .A(n807), .B(b_in[2]), .ZN(n172) );
  INV_X1 U249 ( .A(n172), .ZN(n191) );
  INV_X1 U250 ( .A(n809), .ZN(n171) );
  NAND2_X1 U251 ( .A1(n191), .A2(n334), .ZN(n297) );
  INV_X1 U252 ( .A(n124), .ZN(n174) );
  OR2_X1 U253 ( .A1(n174), .A2(a_in[0]), .ZN(n173) );
  INV_X2 U254 ( .A(n172), .ZN(n372) );
  OAI22_X1 U255 ( .A1(n297), .A2(n174), .B1(n173), .B2(n372), .ZN(n196) );
  NAND2_X1 U256 ( .A1(n191), .A2(n334), .ZN(n374) );
  XNOR2_X1 U257 ( .A(n125), .B(a_in[0]), .ZN(n175) );
  XNOR2_X1 U258 ( .A(n125), .B(a_in[1]), .ZN(n192) );
  OAI22_X1 U259 ( .A1(n374), .A2(n175), .B1(n372), .B2(n192), .ZN(n195) );
  INV_X2 U260 ( .A(n807), .ZN(n797) );
  XNOR2_X1 U261 ( .A(n797), .B(a_in[1]), .ZN(n179) );
  OAI22_X1 U262 ( .A1(n365), .A2(n179), .B1(n176), .B2(n843), .ZN(n178) );
  INV_X1 U263 ( .A(n191), .ZN(n336) );
  AND2_X1 U264 ( .A1(n336), .A2(n131), .ZN(n177) );
  FA_X1 U265 ( .A(n178), .B(f[2]), .CI(n177), .CO(n188), .S(n187) );
  OAI22_X1 U266 ( .A1(n179), .A2(n843), .B1(n365), .B2(a_in[0]), .ZN(n180) );
  NOR2_X1 U267 ( .A1(n187), .A2(n186), .ZN(n614) );
  XNOR2_X1 U268 ( .A(n180), .B(n831), .ZN(n184) );
  INV_X1 U269 ( .A(n797), .ZN(n181) );
  OR2_X1 U270 ( .A1(n131), .A2(n181), .ZN(n182) );
  NAND2_X1 U271 ( .A1(n182), .A2(n365), .ZN(n183) );
  NOR2_X1 U272 ( .A1(n184), .A2(n183), .ZN(n626) );
  AND2_X1 U273 ( .A1(n131), .A2(b_in[0]), .ZN(n624) );
  NAND2_X1 U274 ( .A1(n624), .A2(f[0]), .ZN(n629) );
  NAND2_X1 U275 ( .A1(n184), .A2(n183), .ZN(n627) );
  OAI21_X1 U276 ( .B1(n626), .B2(n629), .A(n627), .ZN(n185) );
  INV_X1 U277 ( .A(n185), .ZN(n618) );
  NAND2_X1 U278 ( .A1(n187), .A2(n186), .ZN(n615) );
  OAI21_X1 U279 ( .B1(n614), .B2(n618), .A(n615), .ZN(n619) );
  AOI21_X1 U280 ( .B1(n621), .B2(n619), .A(n620), .ZN(n613) );
  XNOR2_X1 U281 ( .A(n809), .B(n808), .ZN(n201) );
  INV_X1 U282 ( .A(n490), .ZN(n209) );
  AND2_X1 U283 ( .A1(n209), .A2(n131), .ZN(n205) );
  XNOR2_X1 U284 ( .A(n797), .B(a_in[4]), .ZN(n207) );
  OAI22_X1 U285 ( .A1(n365), .A2(n190), .B1(n207), .B2(n843), .ZN(n204) );
  NAND2_X1 U286 ( .A1(n191), .A2(n334), .ZN(n358) );
  XNOR2_X1 U287 ( .A(n125), .B(a_in[2]), .ZN(n206) );
  OAI22_X1 U288 ( .A1(n358), .A2(n192), .B1(n372), .B2(n206), .ZN(n219) );
  HA_X1 U289 ( .A(n193), .B(f[3]), .CO(n218), .S(n197) );
  XNOR2_X1 U290 ( .A(n217), .B(n194), .ZN(n199) );
  FA_X1 U291 ( .A(n197), .B(n196), .CI(n195), .CO(n198), .S(n189) );
  NOR2_X1 U292 ( .A1(n199), .A2(n198), .ZN(n609) );
  NAND2_X1 U293 ( .A1(n199), .A2(n198), .ZN(n610) );
  OAI21_X1 U294 ( .B1(n613), .B2(n609), .A(n610), .ZN(n608) );
  INV_X1 U295 ( .A(n810), .ZN(n331) );
  XNOR2_X1 U296 ( .A(n331), .B(a_in[0]), .ZN(n203) );
  BUF_X2 U297 ( .A(n201), .Z(n490) );
  INV_X1 U298 ( .A(b_in[4]), .ZN(n200) );
  XNOR2_X2 U299 ( .A(b_in[5]), .B(n200), .ZN(n423) );
  NAND2_X1 U300 ( .A1(n421), .A2(n423), .ZN(n344) );
  XNOR2_X1 U301 ( .A(n331), .B(a_in[1]), .ZN(n234) );
  OR2_X1 U302 ( .A1(n421), .A2(n234), .ZN(n202) );
  OAI21_X1 U303 ( .B1(n344), .B2(n203), .A(n202), .ZN(n236) );
  XNOR2_X1 U304 ( .A(n236), .B(n825), .ZN(n240) );
  FA_X1 U305 ( .A(n205), .B(f[4]), .CI(n204), .CO(n239), .S(n217) );
  XNOR2_X1 U306 ( .A(n240), .B(n239), .ZN(n213) );
  XNOR2_X1 U307 ( .A(n125), .B(a_in[3]), .ZN(n235) );
  OAI22_X1 U308 ( .A1(n374), .A2(n206), .B1(n372), .B2(n235), .ZN(n229) );
  XNOR2_X1 U309 ( .A(n797), .B(a_in[5]), .ZN(n225) );
  OAI22_X1 U310 ( .A1(n365), .A2(n207), .B1(n225), .B2(n843), .ZN(n230) );
  XNOR2_X1 U311 ( .A(n229), .B(n230), .ZN(n212) );
  NAND2_X1 U312 ( .A1(n490), .A2(n423), .ZN(n491) );
  INV_X1 U313 ( .A(n787), .ZN(n211) );
  NOR2_X1 U314 ( .A1(n131), .A2(n211), .ZN(n208) );
  NAND2_X1 U315 ( .A1(n209), .A2(n208), .ZN(n210) );
  OAI21_X1 U316 ( .B1(n491), .B2(n211), .A(n210), .ZN(n231) );
  XNOR2_X1 U317 ( .A(n212), .B(n231), .ZN(n237) );
  XNOR2_X1 U318 ( .A(n213), .B(n237), .ZN(n223) );
  NAND2_X1 U319 ( .A1(n608), .A2(n606), .ZN(n224) );
  NAND2_X1 U320 ( .A1(n223), .A2(n222), .ZN(n605) );
  NAND2_X1 U321 ( .A1(n224), .A2(n605), .ZN(n595) );
  INV_X1 U322 ( .A(n293), .ZN(n294) );
  AND2_X1 U323 ( .A1(a_in[0]), .A2(n294), .ZN(n254) );
  XNOR2_X1 U324 ( .A(n797), .B(a_in[6]), .ZN(n255) );
  OAI22_X1 U325 ( .A1(n365), .A2(n225), .B1(n255), .B2(n843), .ZN(n253) );
  INV_X1 U326 ( .A(n231), .ZN(n227) );
  INV_X1 U327 ( .A(n230), .ZN(n226) );
  NAND2_X1 U328 ( .A1(n227), .A2(n226), .ZN(n228) );
  NAND2_X1 U329 ( .A1(n229), .A2(n228), .ZN(n233) );
  NAND2_X1 U330 ( .A1(n231), .A2(n230), .ZN(n232) );
  NAND2_X1 U331 ( .A1(n233), .A2(n232), .ZN(n261) );
  NAND2_X1 U332 ( .A1(n490), .A2(n423), .ZN(n279) );
  XNOR2_X1 U333 ( .A(n331), .B(a_in[2]), .ZN(n247) );
  OAI22_X1 U334 ( .A1(n279), .A2(n234), .B1(n490), .B2(n247), .ZN(n245) );
  XNOR2_X1 U335 ( .A(n125), .B(a_in[4]), .ZN(n252) );
  OAI22_X1 U336 ( .A1(n297), .A2(n235), .B1(n372), .B2(n252), .ZN(n244) );
  AND2_X1 U337 ( .A1(n236), .A2(f[5]), .ZN(n243) );
  FA_X1 U338 ( .A(n245), .B(n244), .CI(n243), .CO(n286), .S(n260) );
  XNOR2_X1 U339 ( .A(b_in[7]), .B(n811), .ZN(n292) );
  NAND2_X1 U340 ( .A1(n293), .A2(n292), .ZN(n500) );
  OR2_X1 U341 ( .A1(a_in[0]), .A2(n842), .ZN(n246) );
  BUF_X2 U342 ( .A(n293), .Z(n368) );
  OAI22_X1 U343 ( .A1(n500), .A2(n842), .B1(n246), .B2(n368), .ZN(n271) );
  INV_X1 U344 ( .A(n247), .ZN(n249) );
  AND2_X1 U345 ( .A1(n423), .A2(n421), .ZN(n248) );
  NAND2_X1 U346 ( .A1(n249), .A2(n248), .ZN(n251) );
  XNOR2_X1 U347 ( .A(n787), .B(a_in[3]), .ZN(n278) );
  OR2_X1 U348 ( .A1(n278), .A2(n490), .ZN(n250) );
  NAND2_X1 U349 ( .A1(n251), .A2(n250), .ZN(n270) );
  XNOR2_X1 U350 ( .A(n125), .B(a_in[5]), .ZN(n281) );
  OAI22_X1 U351 ( .A1(n374), .A2(n252), .B1(n372), .B2(n281), .ZN(n269) );
  XNOR2_X1 U352 ( .A(n286), .B(n285), .ZN(n259) );
  FA_X1 U353 ( .A(n254), .B(f[6]), .CI(n253), .CO(n274), .S(n262) );
  XNOR2_X1 U354 ( .A(n797), .B(a_in[7]), .ZN(n267) );
  OAI22_X1 U355 ( .A1(n365), .A2(n255), .B1(n267), .B2(n843), .ZN(n273) );
  XNOR2_X1 U356 ( .A(n274), .B(n273), .ZN(n258) );
  NAND2_X1 U357 ( .A1(n293), .A2(n292), .ZN(n370) );
  XNOR2_X1 U358 ( .A(n772), .B(a_in[0]), .ZN(n257) );
  XNOR2_X1 U359 ( .A(b_in[7]), .B(a_in[1]), .ZN(n280) );
  OR2_X1 U360 ( .A1(n368), .A2(n280), .ZN(n256) );
  OAI21_X1 U361 ( .B1(n370), .B2(n257), .A(n256), .ZN(n268) );
  XNOR2_X1 U362 ( .A(n268), .B(n822), .ZN(n272) );
  XNOR2_X1 U363 ( .A(n259), .B(n284), .ZN(n266) );
  FA_X1 U364 ( .A(n262), .B(n261), .CI(n260), .CO(n265), .S(n264) );
  OR2_X2 U365 ( .A1(n266), .A2(n265), .ZN(n597) );
  NAND3_X1 U366 ( .A1(n602), .A2(n595), .A3(n597), .ZN(n593) );
  AND2_X2 U367 ( .A1(n264), .A2(n263), .ZN(n600) );
  NAND2_X1 U368 ( .A1(n600), .A2(n597), .ZN(n592) );
  NAND2_X1 U369 ( .A1(n266), .A2(n265), .ZN(n596) );
  NAND3_X1 U370 ( .A1(n592), .A2(n593), .A3(n596), .ZN(n330) );
  XNOR2_X1 U371 ( .A(n842), .B(n812), .ZN(n298) );
  INV_X1 U372 ( .A(n298), .ZN(n306) );
  AND2_X1 U373 ( .A1(n131), .A2(n306), .ZN(n311) );
  XNOR2_X1 U374 ( .A(b_in[1]), .B(a_in[8]), .ZN(n304) );
  OAI22_X1 U375 ( .A1(n365), .A2(n267), .B1(n304), .B2(n843), .ZN(n310) );
  AND2_X1 U376 ( .A1(n268), .A2(f[7]), .ZN(n290) );
  FA_X1 U377 ( .A(n271), .B(n270), .CI(n269), .CO(n289), .S(n285) );
  XNOR2_X1 U378 ( .A(b_in[5]), .B(a_in[4]), .ZN(n300) );
  OAI22_X1 U379 ( .A1(n279), .A2(n278), .B1(n490), .B2(n300), .ZN(n314) );
  XNOR2_X1 U380 ( .A(n772), .B(a_in[2]), .ZN(n295) );
  OAI22_X1 U381 ( .A1(n500), .A2(n280), .B1(n368), .B2(n295), .ZN(n313) );
  XNOR2_X1 U382 ( .A(n125), .B(a_in[6]), .ZN(n296) );
  OAI22_X1 U383 ( .A1(n297), .A2(n281), .B1(n372), .B2(n296), .ZN(n312) );
  XNOR2_X1 U384 ( .A(n320), .B(n319), .ZN(n282) );
  NOR2_X1 U385 ( .A1(n324), .A2(n323), .ZN(n639) );
  FA_X1 U386 ( .A(n291), .B(n290), .CI(n289), .CO(n461), .S(n318) );
  NAND2_X1 U387 ( .A1(n293), .A2(n292), .ZN(n518) );
  INV_X1 U388 ( .A(n294), .ZN(n519) );
  XNOR2_X1 U389 ( .A(n772), .B(a_in[3]), .ZN(n369) );
  OAI22_X1 U390 ( .A1(n518), .A2(n295), .B1(n519), .B2(n369), .ZN(n395) );
  XNOR2_X1 U391 ( .A(n125), .B(a_in[7]), .ZN(n373) );
  OAI22_X1 U392 ( .A1(n297), .A2(n296), .B1(n372), .B2(n373), .ZN(n394) );
  XNOR2_X1 U393 ( .A(N47), .B(n812), .ZN(n354) );
  XNOR2_X1 U394 ( .A(n842), .B(n812), .ZN(n353) );
  NAND2_X1 U395 ( .A1(n354), .A2(n353), .ZN(n494) );
  XNOR2_X1 U396 ( .A(N47), .B(a_in[0]), .ZN(n299) );
  BUF_X2 U397 ( .A(n298), .Z(n546) );
  XNOR2_X1 U398 ( .A(N47), .B(a_in[1]), .ZN(n377) );
  OAI22_X1 U399 ( .A1(n494), .A2(n299), .B1(n298), .B2(n377), .ZN(n375) );
  XNOR2_X1 U400 ( .A(n375), .B(n826), .ZN(n393) );
  XNOR2_X1 U401 ( .A(n461), .B(n460), .ZN(n316) );
  INV_X1 U402 ( .A(n300), .ZN(n301) );
  NAND3_X1 U403 ( .A1(n423), .A2(n301), .A3(n490), .ZN(n303) );
  XOR2_X1 U404 ( .A(b_in[5]), .B(n806), .Z(n347) );
  OR2_X1 U405 ( .A1(n347), .A2(n421), .ZN(n302) );
  NAND2_X1 U406 ( .A1(n303), .A2(n302), .ZN(n387) );
  XNOR2_X1 U407 ( .A(n797), .B(N46), .ZN(n364) );
  OAI22_X1 U408 ( .A1(n365), .A2(n304), .B1(n364), .B2(n843), .ZN(n385) );
  XNOR2_X1 U409 ( .A(n387), .B(n385), .ZN(n309) );
  NAND2_X1 U410 ( .A1(n306), .A2(n305), .ZN(n308) );
  OR2_X1 U411 ( .A1(n494), .A2(n813), .ZN(n307) );
  XNOR2_X1 U412 ( .A(n309), .B(n386), .ZN(n443) );
  FA_X1 U413 ( .A(n311), .B(f[8]), .CI(n310), .CO(n444), .S(n291) );
  XNOR2_X1 U414 ( .A(n443), .B(n444), .ZN(n315) );
  FA_X1 U415 ( .A(n314), .B(n313), .CI(n312), .CO(n445), .S(n319) );
  XNOR2_X1 U416 ( .A(n315), .B(n445), .ZN(n459) );
  XNOR2_X1 U417 ( .A(n316), .B(n459), .ZN(n326) );
  OR2_X1 U418 ( .A1(n320), .A2(n319), .ZN(n317) );
  NAND2_X1 U419 ( .A1(n320), .A2(n319), .ZN(n321) );
  NOR2_X1 U420 ( .A1(n326), .A2(n325), .ZN(n641) );
  NOR2_X1 U421 ( .A1(n639), .A2(n641), .ZN(n329) );
  NAND2_X1 U422 ( .A1(n324), .A2(n323), .ZN(n638) );
  NOR2_X1 U423 ( .A1(n326), .A2(n325), .ZN(n327) );
  NAND2_X1 U424 ( .A1(n326), .A2(n325), .ZN(n643) );
  OAI21_X1 U425 ( .B1(n638), .B2(n327), .A(n643), .ZN(n328) );
  AOI21_X1 U426 ( .B1(n330), .B2(n329), .A(n328), .ZN(n552) );
  XNOR2_X1 U427 ( .A(n135), .B(a_in[6]), .ZN(n346) );
  XNOR2_X1 U428 ( .A(n331), .B(a_in[7]), .ZN(n343) );
  OR2_X1 U429 ( .A1(n490), .A2(n343), .ZN(n332) );
  OAI21_X1 U430 ( .B1(n491), .B2(n346), .A(n332), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n809), .B(n805), .ZN(n371) );
  INV_X1 U432 ( .A(n371), .ZN(n333) );
  NAND3_X1 U433 ( .A1(n334), .A2(n372), .A3(n333), .ZN(n339) );
  XOR2_X1 U434 ( .A(n124), .B(N46), .Z(n335) );
  NAND2_X1 U435 ( .A1(n336), .A2(n335), .ZN(n338) );
  NAND3_X1 U436 ( .A1(n339), .A2(n338), .A3(f[11]), .ZN(n337) );
  NAND2_X1 U437 ( .A1(n360), .A2(n337), .ZN(n341) );
  NAND2_X1 U438 ( .A1(n339), .A2(n338), .ZN(n361) );
  NAND2_X1 U439 ( .A1(n361), .A2(n816), .ZN(n340) );
  NAND2_X1 U440 ( .A1(n341), .A2(n340), .ZN(n416) );
  XNOR2_X1 U441 ( .A(n135), .B(a_in[8]), .ZN(n420) );
  OR2_X1 U442 ( .A1(n421), .A2(n420), .ZN(n342) );
  OAI21_X1 U443 ( .B1(n344), .B2(n343), .A(n342), .ZN(n427) );
  XNOR2_X1 U444 ( .A(f[11]), .B(f[12]), .ZN(n345) );
  XNOR2_X1 U445 ( .A(n427), .B(n345), .ZN(n414) );
  XNOR2_X1 U446 ( .A(n416), .B(n414), .ZN(n352) );
  INV_X1 U447 ( .A(n813), .ZN(n521) );
  XNOR2_X1 U448 ( .A(n521), .B(a_in[2]), .ZN(n376) );
  XNOR2_X1 U449 ( .A(n521), .B(a_in[3]), .ZN(n355) );
  OAI22_X1 U450 ( .A1(n494), .A2(n376), .B1(n546), .B2(n355), .ZN(n413) );
  XNOR2_X1 U451 ( .A(b_in[7]), .B(a_in[4]), .ZN(n367) );
  XNOR2_X1 U452 ( .A(n772), .B(a_in[5]), .ZN(n356) );
  OAI22_X1 U453 ( .A1(n518), .A2(n367), .B1(n368), .B2(n356), .ZN(n412) );
  OR2_X1 U454 ( .A1(n346), .A2(n421), .ZN(n350) );
  INV_X1 U455 ( .A(n347), .ZN(n348) );
  NAND3_X1 U456 ( .A1(n348), .A2(n423), .A3(n421), .ZN(n349) );
  NAND2_X1 U457 ( .A1(n350), .A2(n349), .ZN(n397) );
  OR2_X1 U458 ( .A1(n397), .A2(f[10]), .ZN(n351) );
  FA_X1 U459 ( .A(n413), .B(n412), .CI(n351), .CO(n417) );
  XNOR2_X1 U460 ( .A(n352), .B(n417), .ZN(n406) );
  NAND2_X1 U461 ( .A1(n354), .A2(n353), .ZN(n545) );
  XNOR2_X1 U462 ( .A(n521), .B(a_in[4]), .ZN(n430) );
  OAI22_X1 U463 ( .A1(n545), .A2(n355), .B1(n546), .B2(n430), .ZN(n433) );
  XNOR2_X1 U464 ( .A(b_in[7]), .B(a_in[6]), .ZN(n425) );
  OAI22_X1 U465 ( .A1(n500), .A2(n356), .B1(n368), .B2(n425), .ZN(n432) );
  XNOR2_X1 U466 ( .A(n125), .B(N46), .ZN(n357) );
  AOI21_X1 U467 ( .B1(n372), .B2(n358), .A(n357), .ZN(n359) );
  INV_X1 U468 ( .A(n359), .ZN(n431) );
  XNOR2_X1 U469 ( .A(n406), .B(n407), .ZN(n381) );
  XNOR2_X1 U470 ( .A(n361), .B(n816), .ZN(n362) );
  XNOR2_X1 U471 ( .A(n363), .B(n362), .ZN(n384) );
  AOI21_X1 U472 ( .B1(n365), .B2(n843), .A(n364), .ZN(n366) );
  INV_X1 U473 ( .A(n366), .ZN(n392) );
  OAI22_X1 U474 ( .A1(n370), .A2(n369), .B1(n368), .B2(n367), .ZN(n391) );
  OAI22_X1 U475 ( .A1(n374), .A2(n373), .B1(n372), .B2(n371), .ZN(n390) );
  XNOR2_X1 U476 ( .A(n397), .B(f[10]), .ZN(n450) );
  AND2_X1 U477 ( .A1(n375), .A2(f[9]), .ZN(n449) );
  NAND2_X1 U478 ( .A1(n450), .A2(n449), .ZN(n380) );
  OAI22_X1 U479 ( .A1(n545), .A2(n377), .B1(n546), .B2(n376), .ZN(n448) );
  NAND2_X1 U480 ( .A1(n450), .A2(n448), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n449), .A2(n448), .ZN(n378) );
  NAND3_X1 U482 ( .A1(n380), .A2(n379), .A3(n378), .ZN(n382) );
  XNOR2_X1 U483 ( .A(n381), .B(n408), .ZN(n469) );
  FA_X1 U484 ( .A(n384), .B(n383), .CI(n382), .CO(n408), .S(n439) );
  FA_X1 U485 ( .A(n395), .B(n394), .CI(n393), .CO(n442) );
  FA_X1 U486 ( .A(n392), .B(n391), .CI(n390), .CO(n383), .S(n453) );
  OAI21_X1 U487 ( .B1(n442), .B2(n441), .A(n453), .ZN(n396) );
  FA_X1 U488 ( .A(n395), .B(n394), .CI(n393), .CO(n401), .S(n460) );
  NAND2_X1 U489 ( .A1(n401), .A2(n441), .ZN(n402) );
  AND2_X1 U490 ( .A1(n396), .A2(n402), .ZN(n399) );
  OR2_X1 U491 ( .A1(n397), .A2(f[10]), .ZN(n411) );
  INV_X1 U492 ( .A(n437), .ZN(n398) );
  NAND2_X1 U493 ( .A1(n399), .A2(n398), .ZN(n400) );
  NAND2_X1 U494 ( .A1(n439), .A2(n400), .ZN(n405) );
  OAI21_X1 U495 ( .B1(n401), .B2(n441), .A(n453), .ZN(n403) );
  NAND2_X1 U496 ( .A1(n403), .A2(n402), .ZN(n438) );
  NAND2_X1 U497 ( .A1(n438), .A2(n437), .ZN(n404) );
  NAND2_X1 U498 ( .A1(n405), .A2(n404), .ZN(n468) );
  NOR2_X1 U499 ( .A1(n469), .A2(n468), .ZN(n571) );
  OAI21_X1 U500 ( .B1(n408), .B2(n407), .A(n406), .ZN(n410) );
  NAND2_X1 U501 ( .A1(n410), .A2(n409), .ZN(n562) );
  FA_X1 U502 ( .A(n413), .B(n412), .CI(n411), .CO(n415), .S(n437) );
  OAI21_X1 U503 ( .B1(n415), .B2(n416), .A(n414), .ZN(n419) );
  NAND2_X1 U504 ( .A1(n416), .A2(n417), .ZN(n418) );
  NAND2_X1 U505 ( .A1(n419), .A2(n418), .ZN(n477) );
  XNOR2_X1 U506 ( .A(n787), .B(N46), .ZN(n489) );
  INV_X1 U507 ( .A(n420), .ZN(n422) );
  NAND3_X1 U508 ( .A1(n423), .A2(n422), .A3(n490), .ZN(n424) );
  OAI21_X1 U509 ( .B1(n490), .B2(n489), .A(n424), .ZN(n488) );
  XNOR2_X1 U510 ( .A(n772), .B(a_in[7]), .ZN(n486) );
  OAI22_X1 U511 ( .A1(n518), .A2(n425), .B1(n519), .B2(n486), .ZN(n487) );
  XNOR2_X1 U512 ( .A(n477), .B(n476), .ZN(n435) );
  NAND2_X1 U513 ( .A1(n816), .A2(n817), .ZN(n426) );
  NAND2_X1 U514 ( .A1(n427), .A2(n426), .ZN(n429) );
  NAND2_X1 U515 ( .A1(f[11]), .A2(f[12]), .ZN(n428) );
  NAND2_X1 U516 ( .A1(n429), .A2(n428), .ZN(n483) );
  XNOR2_X1 U517 ( .A(n521), .B(a_in[5]), .ZN(n493) );
  OAI22_X1 U518 ( .A1(n545), .A2(n430), .B1(n546), .B2(n493), .ZN(n482) );
  FA_X1 U519 ( .A(n433), .B(n432), .CI(n431), .CO(n481), .S(n407) );
  NOR2_X1 U520 ( .A1(n562), .A2(n561), .ZN(n436) );
  NOR2_X1 U521 ( .A1(n571), .A2(n436), .ZN(n472) );
  XNOR2_X1 U522 ( .A(n438), .B(n437), .ZN(n440) );
  XNOR2_X1 U523 ( .A(n440), .B(n439), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n442), .B(n441), .ZN(n454) );
  XOR2_X1 U525 ( .A(n454), .B(n129), .Z(n452) );
  OAI21_X1 U526 ( .B1(n445), .B2(n444), .A(n443), .ZN(n447) );
  NAND2_X1 U527 ( .A1(n447), .A2(n446), .ZN(n456) );
  NAND2_X1 U528 ( .A1(n456), .A2(n455), .ZN(n451) );
  OAI21_X1 U529 ( .B1(n452), .B2(n122), .A(n451), .ZN(n465) );
  NOR2_X1 U530 ( .A1(n466), .A2(n465), .ZN(n554) );
  XNOR2_X1 U531 ( .A(n454), .B(n129), .ZN(n458) );
  XNOR2_X1 U532 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U533 ( .A(n458), .B(n457), .ZN(n590) );
  OAI21_X1 U534 ( .B1(n460), .B2(n461), .A(n459), .ZN(n463) );
  NAND2_X1 U535 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U536 ( .A1(n463), .A2(n462), .ZN(n589) );
  NOR2_X1 U537 ( .A1(n590), .A2(n589), .ZN(n553) );
  NOR2_X1 U538 ( .A1(n554), .A2(n553), .ZN(n464) );
  NAND2_X1 U539 ( .A1(n134), .A2(n464), .ZN(n474) );
  NOR2_X1 U540 ( .A1(n466), .A2(n465), .ZN(n652) );
  NAND2_X1 U541 ( .A1(n590), .A2(n589), .ZN(n467) );
  NAND2_X1 U542 ( .A1(n466), .A2(n465), .ZN(n653) );
  OAI21_X1 U543 ( .B1(n652), .B2(n467), .A(n653), .ZN(n556) );
  NOR2_X1 U544 ( .A1(n562), .A2(n127), .ZN(n470) );
  NAND2_X1 U545 ( .A1(n469), .A2(n468), .ZN(n572) );
  NAND2_X1 U546 ( .A1(n561), .A2(n562), .ZN(n563) );
  OAI21_X1 U547 ( .B1(n470), .B2(n572), .A(n563), .ZN(n471) );
  AOI21_X1 U548 ( .B1(n556), .B2(n472), .A(n471), .ZN(n473) );
  OAI21_X1 U549 ( .B1(n552), .B2(n474), .A(n473), .ZN(n584) );
  INV_X1 U550 ( .A(n584), .ZN(n576) );
  OAI21_X1 U551 ( .B1(n477), .B2(n476), .A(n475), .ZN(n479) );
  NAND2_X1 U552 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U553 ( .A(b_in[7]), .B(a_in[8]), .ZN(n499) );
  OAI22_X1 U554 ( .A1(n500), .A2(n486), .B1(n519), .B2(n499), .ZN(n502) );
  FA_X1 U555 ( .A(n488), .B(n818), .CI(n487), .CO(n503), .S(n476) );
  AOI21_X1 U556 ( .B1(n491), .B2(n490), .A(n489), .ZN(n492) );
  INV_X1 U557 ( .A(n492), .ZN(n505) );
  XNOR2_X1 U558 ( .A(N47), .B(a_in[6]), .ZN(n501) );
  OAI22_X1 U559 ( .A1(n494), .A2(n493), .B1(n546), .B2(n501), .ZN(n504) );
  OR2_X1 U560 ( .A1(n496), .A2(n497), .ZN(n566) );
  INV_X1 U561 ( .A(n566), .ZN(n498) );
  OAI21_X1 U562 ( .B1(n576), .B2(n498), .A(n567), .ZN(n514) );
  XNOR2_X1 U563 ( .A(b_in[7]), .B(N46), .ZN(n517) );
  OAI22_X1 U564 ( .A1(n500), .A2(n499), .B1(n519), .B2(n517), .ZN(n516) );
  XNOR2_X1 U565 ( .A(n521), .B(a_in[7]), .ZN(n522) );
  OAI22_X1 U566 ( .A1(n545), .A2(n501), .B1(n546), .B2(n522), .ZN(n515) );
  FA_X1 U567 ( .A(f[13]), .B(f[14]), .CI(n502), .CO(n524), .S(n509) );
  FA_X1 U568 ( .A(n510), .B(n509), .CI(n508), .CO(n511), .S(n497) );
  NAND2_X1 U569 ( .A1(n512), .A2(n511), .ZN(n533) );
  NAND2_X1 U570 ( .A1(n535), .A2(n533), .ZN(n513) );
  XNOR2_X1 U571 ( .A(n514), .B(n513), .ZN(n719) );
  NAND2_X1 U572 ( .A1(n535), .A2(n566), .ZN(n575) );
  FA_X1 U573 ( .A(n516), .B(n819), .CI(n515), .CO(n530), .S(n525) );
  AOI21_X1 U574 ( .B1(n519), .B2(n518), .A(n517), .ZN(n520) );
  INV_X1 U575 ( .A(n520), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n521), .B(a_in[8]), .ZN(n526) );
  OAI22_X1 U577 ( .A1(n545), .A2(n522), .B1(n546), .B2(n526), .ZN(n527) );
  FA_X1 U578 ( .A(n525), .B(n524), .CI(n523), .CO(n536), .S(n512) );
  NOR2_X1 U579 ( .A1(n537), .A2(n536), .ZN(n577) );
  NOR2_X1 U580 ( .A1(n575), .A2(n577), .ZN(n583) );
  INV_X1 U581 ( .A(n583), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n521), .B(N46), .ZN(n544) );
  OAI22_X1 U583 ( .A1(n545), .A2(n526), .B1(n546), .B2(n544), .ZN(n543) );
  FA_X1 U584 ( .A(f[15]), .B(f[16]), .CI(n527), .CO(n542), .S(n528) );
  FA_X1 U585 ( .A(n530), .B(n529), .CI(n528), .CO(n539), .S(n537) );
  NOR2_X1 U586 ( .A1(n540), .A2(n539), .ZN(n538) );
  NOR2_X1 U587 ( .A1(n531), .A2(n538), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n584), .A2(n532), .ZN(n667) );
  INV_X1 U589 ( .A(n533), .ZN(n534) );
  AOI21_X1 U590 ( .B1(n143), .B2(n535), .A(n534), .ZN(n574) );
  NAND2_X1 U591 ( .A1(n537), .A2(n536), .ZN(n578) );
  OAI21_X1 U592 ( .B1(n574), .B2(n577), .A(n578), .ZN(n582) );
  INV_X1 U593 ( .A(n538), .ZN(n586) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n585) );
  INV_X1 U595 ( .A(n585), .ZN(n541) );
  AOI21_X1 U596 ( .B1(n582), .B2(n586), .A(n541), .ZN(n663) );
  NAND2_X1 U597 ( .A1(n667), .A2(n663), .ZN(n551) );
  FA_X1 U598 ( .A(n543), .B(n820), .CI(n542), .CO(n549), .S(n540) );
  AOI21_X1 U599 ( .B1(n546), .B2(n545), .A(n544), .ZN(n547) );
  INV_X1 U600 ( .A(n547), .ZN(n668) );
  NAND2_X1 U601 ( .A1(n549), .A2(n548), .ZN(n662) );
  NAND2_X1 U602 ( .A1(n661), .A2(n662), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n551), .B(n550), .ZN(n729) );
  NOR2_X1 U604 ( .A1(n719), .A2(n729), .ZN(n660) );
  INV_X1 U605 ( .A(n552), .ZN(n651) );
  NOR2_X1 U606 ( .A1(n554), .A2(n588), .ZN(n570) );
  INV_X1 U607 ( .A(n571), .ZN(n558) );
  AND2_X1 U608 ( .A1(n570), .A2(n558), .ZN(n555) );
  NAND2_X1 U609 ( .A1(n651), .A2(n555), .ZN(n560) );
  AOI21_X1 U610 ( .B1(n569), .B2(n558), .A(n557), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n560), .A2(n559), .ZN(n565) );
  NAND2_X1 U612 ( .A1(n168), .A2(n563), .ZN(n564) );
  XNOR2_X1 U613 ( .A(n565), .B(n564), .ZN(n732) );
  AND2_X1 U614 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U615 ( .A(n576), .B(n568), .ZN(n714) );
  AOI21_X1 U616 ( .B1(n651), .B2(n570), .A(n569), .ZN(n573) );
  XNOR2_X1 U617 ( .A(n573), .B(n169), .ZN(n735) );
  NOR3_X1 U618 ( .A1(n732), .A2(n714), .A3(n735), .ZN(n659) );
  OAI21_X1 U619 ( .B1(n576), .B2(n575), .A(n574), .ZN(n581) );
  INV_X1 U620 ( .A(n577), .ZN(n579) );
  NAND2_X1 U621 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U622 ( .A(n581), .B(n580), .ZN(n726) );
  INV_X1 U623 ( .A(n726), .ZN(n658) );
  AOI21_X1 U624 ( .B1(n584), .B2(n583), .A(n582), .ZN(n587) );
  XNOR2_X1 U625 ( .A(n587), .B(n151), .ZN(n723) );
  INV_X1 U626 ( .A(n588), .ZN(n650) );
  AND2_X1 U627 ( .A1(n590), .A2(n589), .ZN(n649) );
  XNOR2_X1 U628 ( .A(n651), .B(n152), .ZN(n744) );
  INV_X1 U629 ( .A(n639), .ZN(n591) );
  NAND2_X1 U630 ( .A1(n591), .A2(n638), .ZN(n594) );
  AND3_X1 U631 ( .A1(n593), .A2(n592), .A3(n596), .ZN(n640) );
  XNOR2_X1 U632 ( .A(n594), .B(n640), .ZN(n709) );
  BUF_X1 U633 ( .A(n595), .Z(n604) );
  AOI21_X1 U634 ( .B1(n604), .B2(n139), .A(n600), .ZN(n599) );
  NAND2_X1 U635 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U636 ( .A(n599), .B(n598), .Z(n751) );
  INV_X1 U637 ( .A(n600), .ZN(n601) );
  NAND2_X1 U638 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U639 ( .A(n604), .B(n603), .ZN(n754) );
  INV_X1 U640 ( .A(n754), .ZN(n635) );
  NAND2_X1 U641 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U642 ( .A(n137), .B(n607), .ZN(n741) );
  INV_X1 U643 ( .A(n609), .ZN(n611) );
  NAND2_X1 U644 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U645 ( .A(n138), .B(n612), .Z(n757) );
  INV_X1 U646 ( .A(n757), .ZN(n632) );
  INV_X1 U647 ( .A(n614), .ZN(n616) );
  NAND2_X1 U648 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U649 ( .A(n618), .B(n617), .Z(n763) );
  XNOR2_X1 U650 ( .A(n619), .B(n623), .ZN(n760) );
  OR2_X1 U651 ( .A1(n624), .A2(f[0]), .ZN(n625) );
  AND2_X1 U652 ( .A1(n625), .A2(n629), .ZN(n685) );
  INV_X1 U653 ( .A(n626), .ZN(n628) );
  NAND2_X1 U654 ( .A1(n628), .A2(n627), .ZN(n630) );
  XOR2_X1 U655 ( .A(n630), .B(n629), .Z(n766) );
  NOR4_X1 U656 ( .A1(n763), .A2(n760), .A3(n685), .A4(n766), .ZN(n631) );
  NAND2_X1 U657 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U658 ( .A1(n741), .A2(n633), .ZN(n634) );
  NAND2_X1 U659 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U660 ( .A1(n751), .A2(n636), .ZN(n637) );
  AND2_X1 U661 ( .A1(n709), .A2(n637), .ZN(n648) );
  OAI21_X1 U662 ( .B1(n640), .B2(n639), .A(n638), .ZN(n646) );
  INV_X1 U663 ( .A(n642), .ZN(n644) );
  NAND2_X1 U664 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U665 ( .A(n646), .B(n645), .ZN(n748) );
  INV_X1 U666 ( .A(n748), .ZN(n647) );
  NAND3_X1 U667 ( .A1(n744), .A2(n648), .A3(n647), .ZN(n656) );
  AOI21_X1 U668 ( .B1(n651), .B2(n650), .A(n649), .ZN(n655) );
  INV_X1 U669 ( .A(n652), .ZN(n654) );
  XNOR2_X1 U670 ( .A(n655), .B(n147), .ZN(n738) );
  NOR3_X1 U671 ( .A1(n723), .A2(n656), .A3(n738), .ZN(n657) );
  NAND4_X1 U672 ( .A1(n660), .A2(n659), .A3(n658), .A4(n657), .ZN(n684) );
  OAI21_X1 U673 ( .B1(n663), .B2(n666), .A(n662), .ZN(n664) );
  INV_X1 U674 ( .A(n664), .ZN(n665) );
  OAI21_X1 U675 ( .B1(n667), .B2(n666), .A(n665), .ZN(n686) );
  FA_X1 U676 ( .A(f[17]), .B(f[18]), .CI(n668), .CO(n669), .S(n548) );
  XNOR2_X1 U677 ( .A(n686), .B(n146), .ZN(n789) );
  NOR3_X1 U678 ( .A1(n131), .A2(a_in[7]), .A3(a_in[8]), .ZN(n673) );
  NOR2_X1 U679 ( .A1(a_in[5]), .A2(a_in[6]), .ZN(n672) );
  NOR2_X1 U680 ( .A1(a_in[3]), .A2(a_in[4]), .ZN(n671) );
  NOR2_X1 U681 ( .A1(a_in[2]), .A2(a_in[1]), .ZN(n670) );
  NAND4_X1 U682 ( .A1(n673), .A2(n672), .A3(n671), .A4(n670), .ZN(n687) );
  AND2_X1 U683 ( .A1(n687), .A2(N47), .ZN(n681) );
  INV_X1 U684 ( .A(n808), .ZN(n674) );
  NOR3_X1 U685 ( .A1(n132), .A2(b_in[6]), .A3(n674), .ZN(n678) );
  NOR2_X1 U686 ( .A1(b_in[8]), .A2(n778), .ZN(n677) );
  INV_X1 U687 ( .A(n842), .ZN(n772) );
  NOR2_X1 U688 ( .A1(n772), .A2(b_in[0]), .ZN(n676) );
  NOR2_X1 U689 ( .A1(n787), .A2(n171), .ZN(n675) );
  NAND4_X1 U690 ( .A1(n678), .A2(n677), .A3(n676), .A4(n675), .ZN(n679) );
  NAND2_X1 U691 ( .A1(n679), .A2(n813), .ZN(n689) );
  NAND2_X1 U692 ( .A1(n689), .A2(N46), .ZN(n680) );
  OAI211_X1 U693 ( .C1(n681), .C2(N46), .A(N55), .B(n680), .ZN(n682) );
  NOR2_X1 U694 ( .A1(n789), .A2(n682), .ZN(n683) );
  NAND2_X1 U695 ( .A1(n684), .A2(n683), .ZN(n788) );
  NOR2_X1 U696 ( .A1(n814), .A2(reset), .ZN(n844) );
  NAND2_X1 U697 ( .A1(n767), .A2(n685), .ZN(n708) );
  XNOR2_X1 U698 ( .A(n686), .B(n146), .ZN(n705) );
  INV_X1 U699 ( .A(n687), .ZN(n688) );
  OR2_X1 U700 ( .A1(n689), .A2(n688), .ZN(n703) );
  OR2_X1 U701 ( .A1(f[18]), .A2(f[1]), .ZN(n690) );
  NOR3_X1 U702 ( .A1(n690), .A2(f[5]), .A3(f[3]), .ZN(n694) );
  NOR3_X1 U703 ( .A1(f[0]), .A2(f[9]), .A3(f[7]), .ZN(n693) );
  NOR2_X1 U704 ( .A1(f[15]), .A2(f[13]), .ZN(n692) );
  NOR2_X1 U705 ( .A1(f[10]), .A2(f[11]), .ZN(n691) );
  NAND4_X1 U706 ( .A1(n694), .A2(n693), .A3(n692), .A4(n691), .ZN(n701) );
  NOR2_X1 U707 ( .A1(f[16]), .A2(f[14]), .ZN(n698) );
  NOR2_X1 U708 ( .A1(f[12]), .A2(f[8]), .ZN(n697) );
  NOR2_X1 U709 ( .A1(f[6]), .A2(f[4]), .ZN(n696) );
  NOR2_X1 U710 ( .A1(f[17]), .A2(f[2]), .ZN(n695) );
  NAND4_X1 U711 ( .A1(n698), .A2(n697), .A3(n696), .A4(n695), .ZN(n700) );
  AOI21_X1 U712 ( .B1(n813), .B2(N46), .A(N55), .ZN(n699) );
  OAI21_X1 U713 ( .B1(n701), .B2(n700), .A(n699), .ZN(n702) );
  AOI21_X1 U714 ( .B1(n121), .B2(n703), .A(n702), .ZN(n704) );
  OR2_X1 U715 ( .A1(enable_f), .A2(reset), .ZN(n795) );
  NOR2_X1 U716 ( .A1(n795), .A2(n815), .ZN(n706) );
  NOR2_X1 U717 ( .A1(n716), .A2(n706), .ZN(n707) );
  NAND2_X1 U718 ( .A1(n708), .A2(n707), .ZN(n100) );
  NAND2_X1 U719 ( .A1(n133), .A2(n710), .ZN(n713) );
  NOR2_X1 U720 ( .A1(n795), .A2(n830), .ZN(n711) );
  NOR2_X1 U721 ( .A1(n716), .A2(n711), .ZN(n712) );
  NAND2_X1 U722 ( .A1(n713), .A2(n712), .ZN(n92) );
  NAND2_X1 U723 ( .A1(n767), .A2(n714), .ZN(n718) );
  INV_X1 U724 ( .A(n768), .ZN(n716) );
  NOR2_X1 U725 ( .A1(n795), .A2(n827), .ZN(n715) );
  NOR2_X1 U726 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U727 ( .A1(n718), .A2(n717), .ZN(n86) );
  NAND2_X1 U728 ( .A1(n133), .A2(n720), .ZN(n722) );
  NAND2_X1 U729 ( .A1(n722), .A2(n721), .ZN(n85) );
  NAND2_X1 U730 ( .A1(n144), .A2(n723), .ZN(n725) );
  AND2_X1 U731 ( .A1(n768), .A2(n153), .ZN(n724) );
  NAND2_X1 U732 ( .A1(n725), .A2(n724), .ZN(n83) );
  NAND2_X1 U733 ( .A1(n767), .A2(n726), .ZN(n728) );
  AND2_X1 U734 ( .A1(n768), .A2(n154), .ZN(n727) );
  NAND2_X1 U735 ( .A1(n728), .A2(n727), .ZN(n84) );
  NAND2_X1 U736 ( .A1(n133), .A2(n729), .ZN(n731) );
  AND2_X1 U737 ( .A1(n768), .A2(n155), .ZN(n730) );
  NAND2_X1 U738 ( .A1(n731), .A2(n730), .ZN(n82) );
  NAND2_X1 U739 ( .A1(n133), .A2(n732), .ZN(n734) );
  AND2_X1 U740 ( .A1(n768), .A2(n156), .ZN(n733) );
  NAND2_X1 U741 ( .A1(n734), .A2(n733), .ZN(n87) );
  NAND2_X1 U742 ( .A1(n145), .A2(n735), .ZN(n737) );
  AND2_X1 U743 ( .A1(n768), .A2(n157), .ZN(n736) );
  NAND2_X1 U744 ( .A1(n737), .A2(n736), .ZN(n88) );
  NAND2_X1 U745 ( .A1(n145), .A2(n738), .ZN(n740) );
  AND2_X1 U746 ( .A1(n768), .A2(n158), .ZN(n739) );
  NAND2_X1 U747 ( .A1(n740), .A2(n739), .ZN(n89) );
  NAND2_X1 U748 ( .A1(n767), .A2(n741), .ZN(n743) );
  AND2_X1 U749 ( .A1(n768), .A2(n159), .ZN(n742) );
  NAND2_X1 U750 ( .A1(n743), .A2(n742), .ZN(n95) );
  INV_X1 U751 ( .A(n744), .ZN(n745) );
  NAND2_X1 U752 ( .A1(n144), .A2(n745), .ZN(n747) );
  AND2_X1 U753 ( .A1(n768), .A2(n160), .ZN(n746) );
  NAND2_X1 U754 ( .A1(n747), .A2(n746), .ZN(n90) );
  NAND2_X1 U755 ( .A1(n767), .A2(n748), .ZN(n750) );
  AND2_X1 U756 ( .A1(n768), .A2(n161), .ZN(n749) );
  NAND2_X1 U757 ( .A1(n750), .A2(n749), .ZN(n91) );
  NAND2_X1 U758 ( .A1(n145), .A2(n751), .ZN(n753) );
  AND2_X1 U759 ( .A1(n768), .A2(n162), .ZN(n752) );
  NAND2_X1 U760 ( .A1(n753), .A2(n752), .ZN(n93) );
  NAND2_X1 U761 ( .A1(n144), .A2(n754), .ZN(n756) );
  AND2_X1 U762 ( .A1(n768), .A2(n163), .ZN(n755) );
  NAND2_X1 U763 ( .A1(n756), .A2(n755), .ZN(n94) );
  NAND2_X1 U764 ( .A1(n145), .A2(n757), .ZN(n759) );
  AND2_X1 U765 ( .A1(n768), .A2(n164), .ZN(n758) );
  NAND2_X1 U766 ( .A1(n759), .A2(n758), .ZN(n96) );
  NAND2_X1 U767 ( .A1(n144), .A2(n760), .ZN(n762) );
  AND2_X1 U768 ( .A1(n768), .A2(n165), .ZN(n761) );
  NAND2_X1 U769 ( .A1(n762), .A2(n761), .ZN(n97) );
  NAND2_X1 U770 ( .A1(n144), .A2(n763), .ZN(n765) );
  AND2_X1 U771 ( .A1(n768), .A2(n166), .ZN(n764) );
  NAND2_X1 U772 ( .A1(n765), .A2(n764), .ZN(n98) );
  NAND2_X1 U773 ( .A1(n133), .A2(n766), .ZN(n770) );
  AND2_X1 U774 ( .A1(n768), .A2(n167), .ZN(n769) );
  NAND2_X1 U775 ( .A1(n770), .A2(n769), .ZN(n99) );
  INV_X1 U776 ( .A(valid_in), .ZN(n771) );
  NOR2_X2 U777 ( .A1(n771), .A2(reset), .ZN(n800) );
  NOR2_X2 U778 ( .A1(valid_in), .A2(reset), .ZN(n799) );
  AOI22_X1 U779 ( .A1(n800), .A2(b[7]), .B1(n772), .B2(n799), .ZN(n773) );
  INV_X1 U780 ( .A(n773), .ZN(n108) );
  AOI22_X1 U781 ( .A1(n800), .A2(b[3]), .B1(n125), .B2(n799), .ZN(n774) );
  INV_X1 U782 ( .A(n774), .ZN(n104) );
  INV_X1 U783 ( .A(reset), .ZN(n776) );
  INV_X1 U784 ( .A(n800), .ZN(n775) );
  OAI21_X1 U785 ( .B1(n814), .B2(n776), .A(n775), .ZN(n80) );
  AOI22_X1 U786 ( .A1(n800), .A2(b[4]), .B1(n674), .B2(n799), .ZN(n777) );
  INV_X1 U787 ( .A(n777), .ZN(n105) );
  AOI22_X1 U788 ( .A1(n800), .A2(b[2]), .B1(n778), .B2(n799), .ZN(n779) );
  INV_X1 U789 ( .A(n779), .ZN(n103) );
  AOI22_X1 U790 ( .A1(n800), .A2(a[0]), .B1(n131), .B2(n799), .ZN(n780) );
  INV_X1 U791 ( .A(n780), .ZN(n111) );
  AOI22_X1 U792 ( .A1(n800), .A2(a[1]), .B1(a_in[1]), .B2(n799), .ZN(n839) );
  AOI22_X1 U793 ( .A1(n800), .A2(b[6]), .B1(b_in[6]), .B2(n799), .ZN(n781) );
  INV_X1 U794 ( .A(n781), .ZN(n107) );
  AOI22_X1 U795 ( .A1(n800), .A2(a[3]), .B1(a_in[3]), .B2(n799), .ZN(n782) );
  INV_X1 U796 ( .A(n782), .ZN(n114) );
  AOI22_X1 U797 ( .A1(n800), .A2(a[4]), .B1(a_in[4]), .B2(n799), .ZN(n783) );
  INV_X1 U798 ( .A(n783), .ZN(n115) );
  AOI22_X1 U799 ( .A1(n800), .A2(a[5]), .B1(a_in[5]), .B2(n799), .ZN(n838) );
  AOI22_X1 U800 ( .A1(n800), .A2(a[6]), .B1(a_in[6]), .B2(n799), .ZN(n784) );
  INV_X1 U801 ( .A(n784), .ZN(n117) );
  AOI22_X1 U802 ( .A1(n800), .A2(a[2]), .B1(a_in[2]), .B2(n799), .ZN(n785) );
  INV_X1 U803 ( .A(n785), .ZN(n113) );
  AOI22_X1 U804 ( .A1(n800), .A2(a[8]), .B1(a_in[8]), .B2(n799), .ZN(n786) );
  INV_X1 U805 ( .A(n786), .ZN(n119) );
  AOI22_X1 U806 ( .A1(n800), .A2(a[9]), .B1(N46), .B2(n799), .ZN(n836) );
  AOI22_X1 U807 ( .A1(n800), .A2(a[7]), .B1(a_in[7]), .B2(n799), .ZN(n837) );
  AOI22_X1 U808 ( .A1(n800), .A2(b[8]), .B1(b_in[8]), .B2(n799), .ZN(n841) );
  AOI22_X1 U809 ( .A1(n800), .A2(b[5]), .B1(n787), .B2(n799), .ZN(n835) );
  BUF_X1 U810 ( .A(n788), .Z(n792) );
  INV_X1 U811 ( .A(n789), .ZN(n791) );
  INV_X1 U812 ( .A(n844), .ZN(n790) );
  AOI21_X1 U813 ( .B1(n792), .B2(n791), .A(n790), .ZN(n793) );
  NAND2_X1 U814 ( .A1(n141), .A2(n793), .ZN(n794) );
  AOI22_X1 U815 ( .A1(n800), .A2(b[0]), .B1(b_in[0]), .B2(n799), .ZN(n796) );
  INV_X1 U816 ( .A(n796), .ZN(n101) );
  AOI22_X1 U817 ( .A1(n800), .A2(b[1]), .B1(n132), .B2(n799), .ZN(n798) );
  INV_X1 U818 ( .A(n798), .ZN(n102) );
  AOI22_X1 U819 ( .A1(n800), .A2(b[9]), .B1(N47), .B2(n799), .ZN(n840) );
endmodule

