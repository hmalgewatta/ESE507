
module part1_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   enable_f, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527;
  wire   [9:0] a_in;
  wire   [9:0] b_in;

  DFF_X1 enable_f_reg ( .D(n47), .CK(clk), .Q(enable_f), .QN(n525) );
  DFF_X1 \b_in_reg[3]  ( .D(n74), .CK(clk), .Q(b_in[3]), .QN(n527) );
  DFF_X1 valid_out_reg ( .D(n526), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[0]  ( .D(n67), .CK(clk), .Q(f[0]) );
  DFF_X1 \b_in_reg[9]  ( .D(n68), .CK(clk), .Q(b_in[9]), .QN(n522) );
  DFF_X1 \b_in_reg[8]  ( .D(n69), .CK(clk), .Q(b_in[8]) );
  DFF_X1 \b_in_reg[6]  ( .D(n71), .CK(clk), .Q(b_in[6]) );
  DFF_X1 \b_in_reg[5]  ( .D(n72), .CK(clk), .Q(b_in[5]), .QN(n89) );
  DFF_X1 \b_in_reg[4]  ( .D(n73), .CK(clk), .Q(b_in[4]) );
  DFF_X1 \b_in_reg[2]  ( .D(n75), .CK(clk), .Q(b_in[2]), .QN(n524) );
  DFF_X1 \b_in_reg[1]  ( .D(n76), .CK(clk), .Q(b_in[1]), .QN(n523) );
  DFF_X1 \b_in_reg[0]  ( .D(n87), .CK(clk), .Q(b_in[0]), .QN(n521) );
  DFF_X1 \a_in_reg[9]  ( .D(n77), .CK(clk), .Q(a_in[9]) );
  DFF_X1 \a_in_reg[8]  ( .D(n78), .CK(clk), .Q(a_in[8]) );
  DFF_X1 \a_in_reg[7]  ( .D(n79), .CK(clk), .Q(a_in[7]) );
  DFF_X1 \a_in_reg[6]  ( .D(n80), .CK(clk), .Q(a_in[6]) );
  DFF_X1 \a_in_reg[5]  ( .D(n81), .CK(clk), .Q(a_in[5]) );
  DFF_X1 \a_in_reg[4]  ( .D(n82), .CK(clk), .Q(a_in[4]) );
  DFF_X1 \a_in_reg[3]  ( .D(n83), .CK(clk), .Q(a_in[3]) );
  DFF_X1 \a_in_reg[2]  ( .D(n84), .CK(clk), .Q(a_in[2]) );
  DFF_X1 \a_in_reg[1]  ( .D(n85), .CK(clk), .Q(a_in[1]) );
  DFF_X1 \a_in_reg[0]  ( .D(n86), .CK(clk), .Q(a_in[0]) );
  DFF_X1 \f_reg[1]  ( .D(n66), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[2]  ( .D(n65), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(n64), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(n63), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(n62), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[6]  ( .D(n61), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[8]  ( .D(n59), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[7]  ( .D(n60), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[9]  ( .D(n58), .CK(clk), .Q(f[9]) );
  DFF_X1 \f_reg[10]  ( .D(n57), .CK(clk), .Q(f[10]) );
  DFF_X1 \f_reg[11]  ( .D(n56), .CK(clk), .Q(f[11]), .QN(n520) );
  DFF_X1 \f_reg[12]  ( .D(n55), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[13]  ( .D(n54), .CK(clk), .Q(f[13]), .QN(n519) );
  DFF_X1 \f_reg[14]  ( .D(n53), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[17]  ( .D(n50), .CK(clk), .Q(f[17]), .QN(n517) );
  DFF_X1 \f_reg[15]  ( .D(n52), .CK(clk), .Q(f[15]), .QN(n518) );
  DFF_X1 \f_reg[16]  ( .D(n51), .CK(clk), .Q(f[16]) );
  DFF_X1 \f_reg[19]  ( .D(n48), .CK(clk), .Q(f[19]), .QN(n516) );
  DFF_X1 \f_reg[18]  ( .D(n49), .CK(clk), .Q(f[18]) );
  DFF_X2 \b_in_reg[7]  ( .D(n70), .CK(clk), .Q(b_in[7]), .QN(n88) );
  OR2_X1 U91 ( .A1(n237), .A2(n236), .ZN(n247) );
  NAND2_X1 U92 ( .A1(n207), .A2(n206), .ZN(n420) );
  OR2_X1 U93 ( .A1(n306), .A2(n305), .ZN(n357) );
  NAND2_X1 U94 ( .A1(n169), .A2(n149), .ZN(n399) );
  NAND2_X1 U95 ( .A1(n263), .A2(n488), .ZN(n487) );
  NAND2_X1 U96 ( .A1(n306), .A2(n305), .ZN(n90) );
  XNOR2_X1 U97 ( .A(b_in[3]), .B(b_in[4]), .ZN(n149) );
  INV_X1 U98 ( .A(reset), .ZN(n92) );
  AND2_X1 U99 ( .A1(enable_f), .A2(n92), .ZN(n526) );
  AND2_X1 U100 ( .A1(valid_in), .A2(n92), .ZN(n514) );
  INV_X1 U101 ( .A(n514), .ZN(n91) );
  OAI21_X1 U102 ( .B1(n525), .B2(n92), .A(n91), .ZN(n47) );
  AND2_X1 U103 ( .A1(a_in[0]), .A2(b_in[0]), .ZN(n93) );
  OR2_X1 U104 ( .A1(n93), .A2(f[0]), .ZN(n94) );
  NAND2_X1 U105 ( .A1(n93), .A2(f[0]), .ZN(n132) );
  AND2_X1 U106 ( .A1(n94), .A2(n132), .ZN(n95) );
  NOR2_X2 U107 ( .A1(enable_f), .A2(reset), .ZN(n509) );
  AOI22_X1 U108 ( .A1(n95), .A2(n526), .B1(n509), .B2(f[0]), .ZN(n96) );
  INV_X1 U109 ( .A(n96), .ZN(n67) );
  NOR2_X2 U110 ( .A1(valid_in), .A2(reset), .ZN(n513) );
  AOI22_X1 U111 ( .A1(n514), .A2(a[9]), .B1(n513), .B2(a_in[9]), .ZN(n97) );
  INV_X1 U112 ( .A(n97), .ZN(n77) );
  AOI22_X1 U113 ( .A1(n514), .A2(a[8]), .B1(n513), .B2(a_in[8]), .ZN(n98) );
  INV_X1 U114 ( .A(n98), .ZN(n78) );
  AOI22_X1 U115 ( .A1(n514), .A2(b[0]), .B1(n513), .B2(b_in[0]), .ZN(n99) );
  INV_X1 U116 ( .A(n99), .ZN(n87) );
  AOI22_X1 U117 ( .A1(n514), .A2(a[7]), .B1(n513), .B2(a_in[7]), .ZN(n100) );
  INV_X1 U118 ( .A(n100), .ZN(n79) );
  AOI22_X1 U119 ( .A1(n514), .A2(a[6]), .B1(n513), .B2(a_in[6]), .ZN(n101) );
  INV_X1 U120 ( .A(n101), .ZN(n80) );
  AOI22_X1 U121 ( .A1(n514), .A2(a[5]), .B1(n513), .B2(a_in[5]), .ZN(n102) );
  INV_X1 U122 ( .A(n102), .ZN(n81) );
  AOI22_X1 U123 ( .A1(n514), .A2(a[4]), .B1(n513), .B2(a_in[4]), .ZN(n103) );
  INV_X1 U124 ( .A(n103), .ZN(n82) );
  AOI22_X1 U125 ( .A1(n514), .A2(a[0]), .B1(n513), .B2(a_in[0]), .ZN(n104) );
  INV_X1 U126 ( .A(n104), .ZN(n86) );
  AOI22_X1 U127 ( .A1(n514), .A2(a[3]), .B1(n513), .B2(a_in[3]), .ZN(n105) );
  INV_X1 U128 ( .A(n105), .ZN(n83) );
  AOI22_X1 U129 ( .A1(n514), .A2(a[2]), .B1(n513), .B2(a_in[2]), .ZN(n106) );
  INV_X1 U130 ( .A(n106), .ZN(n84) );
  AOI22_X1 U131 ( .A1(n514), .A2(a[1]), .B1(n513), .B2(a_in[1]), .ZN(n107) );
  INV_X1 U132 ( .A(n107), .ZN(n85) );
  AOI22_X1 U133 ( .A1(n514), .A2(b[8]), .B1(n513), .B2(b_in[8]), .ZN(n108) );
  INV_X1 U134 ( .A(n108), .ZN(n69) );
  AOI22_X1 U135 ( .A1(n514), .A2(b[6]), .B1(n513), .B2(b_in[6]), .ZN(n109) );
  INV_X1 U136 ( .A(n109), .ZN(n71) );
  AOI22_X1 U137 ( .A1(n514), .A2(b[4]), .B1(n513), .B2(b_in[4]), .ZN(n110) );
  INV_X1 U138 ( .A(n110), .ZN(n73) );
  AOI22_X1 U139 ( .A1(n514), .A2(b[2]), .B1(n513), .B2(b_in[2]), .ZN(n111) );
  INV_X1 U140 ( .A(n111), .ZN(n75) );
  NAND2_X1 U141 ( .A1(b_in[1]), .A2(n521), .ZN(n294) );
  XNOR2_X1 U142 ( .A(b_in[1]), .B(a_in[1]), .ZN(n125) );
  OAI22_X1 U143 ( .A1(n294), .A2(a_in[0]), .B1(n125), .B2(n521), .ZN(n130) );
  OR2_X1 U144 ( .A1(a_in[0]), .A2(n523), .ZN(n112) );
  NAND2_X1 U145 ( .A1(n112), .A2(n294), .ZN(n113) );
  NOR2_X1 U146 ( .A1(n114), .A2(n113), .ZN(n133) );
  INV_X1 U147 ( .A(n133), .ZN(n115) );
  NAND2_X1 U148 ( .A1(n114), .A2(n113), .ZN(n131) );
  NAND2_X1 U149 ( .A1(n115), .A2(n131), .ZN(n116) );
  XOR2_X1 U150 ( .A(n116), .B(n132), .Z(n117) );
  AOI22_X1 U151 ( .A1(n117), .A2(n526), .B1(n509), .B2(f[1]), .ZN(n118) );
  INV_X1 U152 ( .A(n118), .ZN(n66) );
  XNOR2_X1 U153 ( .A(b_in[2]), .B(b_in[1]), .ZN(n120) );
  XNOR2_X1 U154 ( .A(b_in[3]), .B(n524), .ZN(n119) );
  NAND2_X1 U155 ( .A1(n120), .A2(n119), .ZN(n338) );
  OR2_X1 U156 ( .A1(a_in[0]), .A2(n527), .ZN(n121) );
  BUF_X1 U157 ( .A(n120), .Z(n317) );
  OAI22_X1 U158 ( .A1(n338), .A2(n527), .B1(n121), .B2(n317), .ZN(n153) );
  XNOR2_X1 U159 ( .A(b_in[3]), .B(a_in[0]), .ZN(n122) );
  XNOR2_X1 U160 ( .A(b_in[3]), .B(a_in[1]), .ZN(n148) );
  OAI22_X1 U161 ( .A1(n338), .A2(n122), .B1(n317), .B2(n148), .ZN(n152) );
  XNOR2_X1 U162 ( .A(b_in[1]), .B(a_in[2]), .ZN(n124) );
  XNOR2_X1 U163 ( .A(b_in[1]), .B(a_in[3]), .ZN(n150) );
  OAI22_X1 U164 ( .A1(n294), .A2(n124), .B1(n150), .B2(n521), .ZN(n147) );
  INV_X1 U165 ( .A(n317), .ZN(n123) );
  AND2_X1 U166 ( .A1(a_in[0]), .A2(n123), .ZN(n129) );
  OAI22_X1 U167 ( .A1(n294), .A2(n125), .B1(n124), .B2(n521), .ZN(n128) );
  OR2_X1 U168 ( .A1(n127), .A2(n126), .ZN(n160) );
  NAND2_X1 U169 ( .A1(n127), .A2(n126), .ZN(n157) );
  NAND2_X1 U170 ( .A1(n160), .A2(n157), .ZN(n137) );
  FA_X1 U171 ( .A(n129), .B(f[2]), .CI(n128), .CO(n126), .S(n136) );
  HA_X1 U172 ( .A(n130), .B(f[1]), .CO(n135), .S(n114) );
  NOR2_X1 U173 ( .A1(n136), .A2(n135), .ZN(n140) );
  OAI21_X1 U174 ( .B1(n133), .B2(n132), .A(n131), .ZN(n134) );
  INV_X1 U175 ( .A(n134), .ZN(n143) );
  NAND2_X1 U176 ( .A1(n136), .A2(n135), .ZN(n141) );
  OAI21_X1 U177 ( .B1(n140), .B2(n143), .A(n141), .ZN(n159) );
  XNOR2_X1 U178 ( .A(n137), .B(n159), .ZN(n138) );
  AOI22_X1 U179 ( .A1(n138), .A2(n526), .B1(n509), .B2(f[3]), .ZN(n139) );
  INV_X1 U180 ( .A(n139), .ZN(n64) );
  INV_X1 U181 ( .A(n140), .ZN(n142) );
  NAND2_X1 U182 ( .A1(n142), .A2(n141), .ZN(n144) );
  XOR2_X1 U183 ( .A(n144), .B(n143), .Z(n145) );
  AOI22_X1 U184 ( .A1(n145), .A2(n526), .B1(n509), .B2(f[2]), .ZN(n146) );
  INV_X1 U185 ( .A(n146), .ZN(n65) );
  HA_X1 U186 ( .A(n147), .B(f[3]), .CO(n177), .S(n151) );
  XNOR2_X1 U187 ( .A(b_in[3]), .B(a_in[2]), .ZN(n174) );
  OAI22_X1 U188 ( .A1(n338), .A2(n148), .B1(n120), .B2(n174), .ZN(n176) );
  INV_X1 U189 ( .A(n149), .ZN(n170) );
  AND2_X1 U190 ( .A1(a_in[0]), .A2(n170), .ZN(n168) );
  XNOR2_X1 U191 ( .A(b_in[1]), .B(a_in[4]), .ZN(n173) );
  OAI22_X1 U192 ( .A1(n294), .A2(n150), .B1(n173), .B2(n521), .ZN(n167) );
  FA_X1 U193 ( .A(n153), .B(n152), .CI(n151), .CO(n154), .S(n127) );
  NOR2_X1 U194 ( .A1(n155), .A2(n154), .ZN(n166) );
  INV_X1 U195 ( .A(n166), .ZN(n156) );
  NAND2_X1 U196 ( .A1(n155), .A2(n154), .ZN(n164) );
  NAND2_X1 U197 ( .A1(n156), .A2(n164), .ZN(n161) );
  INV_X1 U198 ( .A(n157), .ZN(n158) );
  AOI21_X1 U199 ( .B1(n160), .B2(n159), .A(n158), .ZN(n165) );
  XOR2_X1 U200 ( .A(n161), .B(n165), .Z(n162) );
  AOI22_X1 U201 ( .A1(n162), .A2(n526), .B1(n509), .B2(f[4]), .ZN(n163) );
  INV_X1 U202 ( .A(n163), .ZN(n63) );
  OAI21_X1 U203 ( .B1(n166), .B2(n165), .A(n164), .ZN(n186) );
  FA_X1 U204 ( .A(n168), .B(f[4]), .CI(n167), .CO(n196), .S(n175) );
  XOR2_X1 U205 ( .A(b_in[4]), .B(b_in[5]), .Z(n169) );
  BUF_X1 U206 ( .A(b_in[5]), .Z(n378) );
  XNOR2_X1 U207 ( .A(n378), .B(a_in[0]), .ZN(n171) );
  INV_X1 U208 ( .A(n170), .ZN(n400) );
  XNOR2_X1 U209 ( .A(n378), .B(a_in[1]), .ZN(n191) );
  OAI22_X1 U210 ( .A1(n399), .A2(n171), .B1(n400), .B2(n191), .ZN(n193) );
  OR2_X1 U211 ( .A1(a_in[0]), .A2(n89), .ZN(n172) );
  OAI22_X1 U212 ( .A1(n399), .A2(n89), .B1(n172), .B2(n400), .ZN(n190) );
  XNOR2_X1 U213 ( .A(b_in[1]), .B(a_in[5]), .ZN(n187) );
  OAI22_X1 U214 ( .A1(n294), .A2(n173), .B1(n187), .B2(n521), .ZN(n189) );
  XNOR2_X1 U215 ( .A(b_in[3]), .B(a_in[3]), .ZN(n192) );
  OAI22_X1 U216 ( .A1(n338), .A2(n174), .B1(n120), .B2(n192), .ZN(n188) );
  FA_X1 U217 ( .A(n177), .B(n176), .CI(n175), .CO(n178), .S(n155) );
  OR2_X1 U218 ( .A1(n179), .A2(n178), .ZN(n185) );
  NAND2_X1 U219 ( .A1(n179), .A2(n178), .ZN(n183) );
  NAND2_X1 U220 ( .A1(n185), .A2(n183), .ZN(n180) );
  XNOR2_X1 U221 ( .A(n186), .B(n180), .ZN(n181) );
  AOI22_X1 U222 ( .A1(n181), .A2(n526), .B1(n509), .B2(f[5]), .ZN(n182) );
  INV_X1 U223 ( .A(n182), .ZN(n62) );
  INV_X1 U224 ( .A(n183), .ZN(n184) );
  AOI21_X1 U225 ( .B1(n186), .B2(n185), .A(n184), .ZN(n239) );
  INV_X1 U226 ( .A(n239), .ZN(n246) );
  XOR2_X1 U227 ( .A(b_in[6]), .B(b_in[5]), .Z(n208) );
  AND2_X1 U228 ( .A1(a_in[0]), .A2(n208), .ZN(n204) );
  XNOR2_X1 U229 ( .A(b_in[1]), .B(a_in[6]), .ZN(n205) );
  OAI22_X1 U230 ( .A1(n294), .A2(n187), .B1(n205), .B2(n521), .ZN(n203) );
  FA_X1 U231 ( .A(n190), .B(n189), .CI(n188), .CO(n234), .S(n194) );
  XNOR2_X1 U232 ( .A(n378), .B(a_in[2]), .ZN(n214) );
  OAI22_X1 U233 ( .A1(n399), .A2(n191), .B1(n400), .B2(n214), .ZN(n224) );
  XNOR2_X1 U234 ( .A(b_in[3]), .B(a_in[4]), .ZN(n212) );
  OAI22_X1 U235 ( .A1(n338), .A2(n192), .B1(n120), .B2(n212), .ZN(n223) );
  HA_X1 U236 ( .A(n193), .B(f[5]), .CO(n222), .S(n195) );
  FA_X1 U237 ( .A(n196), .B(n195), .CI(n194), .CO(n197), .S(n179) );
  OR2_X1 U238 ( .A1(n198), .A2(n197), .ZN(n245) );
  AND2_X1 U239 ( .A1(n198), .A2(n197), .ZN(n244) );
  INV_X1 U240 ( .A(n244), .ZN(n199) );
  NAND2_X1 U241 ( .A1(n245), .A2(n199), .ZN(n200) );
  XNOR2_X1 U242 ( .A(n246), .B(n200), .ZN(n201) );
  AOI22_X1 U243 ( .A1(n201), .A2(n526), .B1(n509), .B2(f[6]), .ZN(n202) );
  INV_X1 U244 ( .A(n202), .ZN(n61) );
  FA_X1 U245 ( .A(n204), .B(f[6]), .CI(n203), .CO(n227), .S(n235) );
  XNOR2_X1 U246 ( .A(b_in[1]), .B(a_in[7]), .ZN(n218) );
  OAI22_X1 U247 ( .A1(n294), .A2(n205), .B1(n218), .B2(n521), .ZN(n226) );
  INV_X1 U248 ( .A(n208), .ZN(n207) );
  XOR2_X1 U249 ( .A(b_in[6]), .B(b_in[7]), .Z(n206) );
  XNOR2_X1 U250 ( .A(b_in[7]), .B(a_in[0]), .ZN(n209) );
  INV_X1 U251 ( .A(n208), .ZN(n421) );
  XNOR2_X1 U252 ( .A(b_in[7]), .B(a_in[1]), .ZN(n210) );
  OAI22_X1 U253 ( .A1(n420), .A2(n209), .B1(n421), .B2(n210), .ZN(n216) );
  XNOR2_X1 U254 ( .A(b_in[7]), .B(a_in[2]), .ZN(n270) );
  OAI22_X1 U255 ( .A1(n420), .A2(n210), .B1(n421), .B2(n270), .ZN(n267) );
  XNOR2_X1 U256 ( .A(b_in[3]), .B(a_in[5]), .ZN(n211) );
  XNOR2_X1 U257 ( .A(b_in[3]), .B(a_in[6]), .ZN(n262) );
  OAI22_X1 U258 ( .A1(n338), .A2(n211), .B1(n120), .B2(n262), .ZN(n266) );
  XNOR2_X1 U259 ( .A(n378), .B(a_in[3]), .ZN(n213) );
  XNOR2_X1 U260 ( .A(n378), .B(a_in[4]), .ZN(n261) );
  OAI22_X1 U261 ( .A1(n399), .A2(n213), .B1(n400), .B2(n261), .ZN(n265) );
  OAI22_X1 U262 ( .A1(n338), .A2(n212), .B1(n317), .B2(n211), .ZN(n221) );
  OAI22_X1 U263 ( .A1(n399), .A2(n214), .B1(n400), .B2(n213), .ZN(n220) );
  OR2_X1 U264 ( .A1(a_in[0]), .A2(n88), .ZN(n215) );
  OAI22_X1 U265 ( .A1(n420), .A2(n88), .B1(n215), .B2(n421), .ZN(n219) );
  HA_X1 U266 ( .A(n216), .B(f[7]), .CO(n259), .S(n225) );
  XNOR2_X2 U267 ( .A(b_in[8]), .B(b_in[7]), .ZN(n488) );
  INV_X1 U268 ( .A(n488), .ZN(n217) );
  AND2_X1 U269 ( .A1(a_in[0]), .A2(n217), .ZN(n269) );
  XNOR2_X1 U270 ( .A(b_in[1]), .B(a_in[8]), .ZN(n272) );
  OAI22_X1 U271 ( .A1(n294), .A2(n218), .B1(n272), .B2(n521), .ZN(n268) );
  FA_X1 U272 ( .A(n221), .B(n220), .CI(n219), .CO(n260), .S(n232) );
  FA_X1 U273 ( .A(n224), .B(n223), .CI(n222), .CO(n231), .S(n233) );
  FA_X1 U274 ( .A(n227), .B(n226), .CI(n225), .CO(n275), .S(n230) );
  OR2_X1 U275 ( .A1(n229), .A2(n228), .ZN(n256) );
  NAND2_X1 U276 ( .A1(n229), .A2(n228), .ZN(n254) );
  NAND2_X1 U277 ( .A1(n256), .A2(n254), .ZN(n241) );
  FA_X1 U278 ( .A(n232), .B(n231), .CI(n230), .CO(n228), .S(n237) );
  FA_X1 U279 ( .A(n235), .B(n234), .CI(n233), .CO(n236), .S(n198) );
  NAND2_X1 U280 ( .A1(n247), .A2(n245), .ZN(n240) );
  AND2_X1 U281 ( .A1(n237), .A2(n236), .ZN(n248) );
  AOI21_X1 U282 ( .B1(n247), .B2(n244), .A(n248), .ZN(n238) );
  OAI21_X1 U283 ( .B1(n240), .B2(n239), .A(n238), .ZN(n257) );
  XNOR2_X1 U284 ( .A(n241), .B(n257), .ZN(n242) );
  AOI22_X1 U285 ( .A1(n242), .A2(n526), .B1(n509), .B2(f[8]), .ZN(n243) );
  INV_X1 U286 ( .A(n243), .ZN(n59) );
  AOI21_X1 U287 ( .B1(n246), .B2(n245), .A(n244), .ZN(n251) );
  INV_X1 U288 ( .A(n248), .ZN(n249) );
  NAND2_X1 U289 ( .A1(n247), .A2(n249), .ZN(n250) );
  XOR2_X1 U290 ( .A(n251), .B(n250), .Z(n252) );
  AOI22_X1 U291 ( .A1(n252), .A2(n526), .B1(n509), .B2(f[7]), .ZN(n253) );
  INV_X1 U292 ( .A(n253), .ZN(n60) );
  INV_X1 U293 ( .A(n254), .ZN(n255) );
  AOI21_X1 U294 ( .B1(n257), .B2(n256), .A(n255), .ZN(n284) );
  FA_X1 U295 ( .A(n260), .B(n259), .CI(n258), .CO(n304), .S(n273) );
  XNOR2_X1 U296 ( .A(n378), .B(a_in[5]), .ZN(n292) );
  OAI22_X1 U297 ( .A1(n399), .A2(n261), .B1(n400), .B2(n292), .ZN(n301) );
  XNOR2_X1 U298 ( .A(b_in[3]), .B(a_in[7]), .ZN(n291) );
  OAI22_X1 U299 ( .A1(n338), .A2(n262), .B1(n317), .B2(n291), .ZN(n300) );
  XOR2_X1 U300 ( .A(b_in[8]), .B(b_in[9]), .Z(n263) );
  OR2_X1 U301 ( .A1(a_in[0]), .A2(n522), .ZN(n264) );
  OAI22_X1 U302 ( .A1(n487), .A2(n522), .B1(n264), .B2(n488), .ZN(n288) );
  FA_X1 U303 ( .A(n267), .B(n266), .CI(n265), .CO(n287), .S(n274) );
  FA_X1 U304 ( .A(n269), .B(f[8]), .CI(n268), .CO(n286), .S(n258) );
  XNOR2_X1 U305 ( .A(b_in[7]), .B(a_in[3]), .ZN(n289) );
  OAI22_X1 U306 ( .A1(n420), .A2(n270), .B1(n421), .B2(n289), .ZN(n298) );
  XNOR2_X1 U307 ( .A(b_in[9]), .B(a_in[0]), .ZN(n271) );
  XNOR2_X1 U308 ( .A(b_in[9]), .B(a_in[1]), .ZN(n290) );
  OAI22_X1 U309 ( .A1(n487), .A2(n271), .B1(n488), .B2(n290), .ZN(n297) );
  XNOR2_X1 U310 ( .A(b_in[1]), .B(a_in[9]), .ZN(n293) );
  OAI22_X1 U311 ( .A1(n294), .A2(n272), .B1(n293), .B2(n521), .ZN(n296) );
  FA_X1 U312 ( .A(n275), .B(n274), .CI(n273), .CO(n276), .S(n229) );
  NOR2_X1 U313 ( .A1(n277), .A2(n276), .ZN(n283) );
  INV_X1 U314 ( .A(n283), .ZN(n278) );
  NAND2_X1 U315 ( .A1(n277), .A2(n276), .ZN(n282) );
  NAND2_X1 U316 ( .A1(n278), .A2(n282), .ZN(n279) );
  XOR2_X1 U317 ( .A(n284), .B(n279), .Z(n280) );
  AOI22_X1 U318 ( .A1(n280), .A2(n526), .B1(n509), .B2(f[9]), .ZN(n281) );
  INV_X1 U319 ( .A(n281), .ZN(n58) );
  OAI21_X1 U320 ( .B1(n284), .B2(n283), .A(n282), .ZN(n367) );
  FA_X1 U321 ( .A(n287), .B(n286), .CI(n285), .CO(n327), .S(n302) );
  HA_X1 U322 ( .A(n288), .B(f[9]), .CO(n324), .S(n299) );
  XNOR2_X1 U323 ( .A(b_in[7]), .B(a_in[4]), .ZN(n313) );
  OAI22_X1 U324 ( .A1(n420), .A2(n289), .B1(n421), .B2(n313), .ZN(n323) );
  XNOR2_X1 U325 ( .A(b_in[9]), .B(a_in[2]), .ZN(n316) );
  OAI22_X1 U326 ( .A1(n487), .A2(n290), .B1(n316), .B2(n488), .ZN(n315) );
  XNOR2_X1 U327 ( .A(n315), .B(f[10]), .ZN(n322) );
  XNOR2_X1 U328 ( .A(b_in[3]), .B(a_in[8]), .ZN(n318) );
  OAI22_X1 U329 ( .A1(n338), .A2(n291), .B1(n317), .B2(n318), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n378), .B(a_in[6]), .ZN(n314) );
  OAI22_X1 U331 ( .A1(n399), .A2(n292), .B1(n400), .B2(n314), .ZN(n320) );
  AOI21_X1 U332 ( .B1(n294), .B2(n521), .A(n293), .ZN(n295) );
  INV_X1 U333 ( .A(n295), .ZN(n319) );
  FA_X1 U334 ( .A(n298), .B(n297), .CI(n296), .CO(n311), .S(n285) );
  FA_X1 U335 ( .A(n301), .B(n300), .CI(n299), .CO(n310), .S(n303) );
  FA_X1 U336 ( .A(n304), .B(n303), .CI(n302), .CO(n305), .S(n277) );
  NAND2_X1 U337 ( .A1(n357), .A2(n90), .ZN(n307) );
  XNOR2_X1 U338 ( .A(n367), .B(n307), .ZN(n308) );
  AOI22_X1 U339 ( .A1(n308), .A2(n526), .B1(n509), .B2(f[10]), .ZN(n309) );
  INV_X1 U340 ( .A(n309), .ZN(n57) );
  FA_X1 U341 ( .A(n312), .B(n311), .CI(n310), .CO(n350), .S(n325) );
  XNOR2_X1 U342 ( .A(b_in[7]), .B(a_in[5]), .ZN(n336) );
  OAI22_X1 U343 ( .A1(n420), .A2(n313), .B1(n421), .B2(n336), .ZN(n344) );
  XNOR2_X1 U344 ( .A(n378), .B(a_in[7]), .ZN(n337) );
  OAI22_X1 U345 ( .A1(n399), .A2(n314), .B1(n400), .B2(n337), .ZN(n343) );
  OR2_X1 U346 ( .A1(n315), .A2(f[10]), .ZN(n342) );
  XNOR2_X1 U347 ( .A(b_in[9]), .B(a_in[3]), .ZN(n347) );
  OAI22_X1 U348 ( .A1(n487), .A2(n316), .B1(n488), .B2(n347), .ZN(n346) );
  XNOR2_X1 U349 ( .A(b_in[3]), .B(a_in[9]), .ZN(n339) );
  OAI22_X1 U350 ( .A1(n338), .A2(n318), .B1(n317), .B2(n339), .ZN(n345) );
  FA_X1 U351 ( .A(n321), .B(n320), .CI(n319), .CO(n334), .S(n312) );
  FA_X1 U352 ( .A(n324), .B(n323), .CI(n322), .CO(n333), .S(n326) );
  FA_X1 U353 ( .A(n327), .B(n326), .CI(n325), .CO(n328), .S(n306) );
  NAND2_X1 U354 ( .A1(n329), .A2(n328), .ZN(n359) );
  NAND2_X1 U355 ( .A1(n90), .A2(n359), .ZN(n365) );
  OR2_X1 U356 ( .A1(n329), .A2(n328), .ZN(n360) );
  INV_X1 U357 ( .A(n360), .ZN(n331) );
  INV_X1 U358 ( .A(n357), .ZN(n330) );
  OAI21_X1 U359 ( .B1(n331), .B2(n330), .A(n359), .ZN(n371) );
  OAI21_X1 U360 ( .B1(n367), .B2(n365), .A(n371), .ZN(n332) );
  INV_X1 U361 ( .A(n332), .ZN(n354) );
  FA_X1 U362 ( .A(n335), .B(n334), .CI(n333), .CO(n387), .S(n348) );
  XNOR2_X1 U363 ( .A(b_in[7]), .B(a_in[6]), .ZN(n381) );
  OAI22_X1 U364 ( .A1(n420), .A2(n336), .B1(n421), .B2(n381), .ZN(n384) );
  XNOR2_X1 U365 ( .A(n378), .B(a_in[8]), .ZN(n379) );
  OAI22_X1 U366 ( .A1(n399), .A2(n337), .B1(n400), .B2(n379), .ZN(n383) );
  NAND2_X1 U367 ( .A1(n338), .A2(n120), .ZN(n341) );
  INV_X1 U368 ( .A(n339), .ZN(n340) );
  NAND2_X1 U369 ( .A1(n341), .A2(n340), .ZN(n382) );
  FA_X1 U370 ( .A(n344), .B(n343), .CI(n342), .CO(n376), .S(n349) );
  FA_X1 U371 ( .A(n346), .B(n520), .CI(n345), .CO(n375), .S(n335) );
  XNOR2_X1 U372 ( .A(b_in[9]), .B(a_in[4]), .ZN(n377) );
  OAI22_X1 U373 ( .A1(n487), .A2(n347), .B1(n488), .B2(n377), .ZN(n380) );
  FA_X1 U374 ( .A(n350), .B(n349), .CI(n348), .CO(n351), .S(n329) );
  OR2_X1 U375 ( .A1(n352), .A2(n351), .ZN(n370) );
  NAND2_X1 U376 ( .A1(n352), .A2(n351), .ZN(n372) );
  NAND2_X1 U377 ( .A1(n370), .A2(n372), .ZN(n353) );
  XNOR2_X1 U378 ( .A(n354), .B(n353), .ZN(n355) );
  AOI22_X1 U379 ( .A1(n355), .A2(n526), .B1(n509), .B2(f[12]), .ZN(n356) );
  INV_X1 U380 ( .A(n356), .ZN(n55) );
  NAND2_X1 U381 ( .A1(n367), .A2(n357), .ZN(n358) );
  NAND2_X1 U382 ( .A1(n358), .A2(n90), .ZN(n362) );
  NAND2_X1 U383 ( .A1(n360), .A2(n359), .ZN(n361) );
  XNOR2_X1 U384 ( .A(n362), .B(n361), .ZN(n363) );
  AOI22_X1 U385 ( .A1(n363), .A2(n526), .B1(n509), .B2(f[11]), .ZN(n364) );
  INV_X1 U386 ( .A(n364), .ZN(n56) );
  INV_X1 U387 ( .A(n372), .ZN(n366) );
  NOR2_X1 U388 ( .A1(n366), .A2(n365), .ZN(n369) );
  INV_X1 U389 ( .A(n367), .ZN(n368) );
  NAND2_X1 U390 ( .A1(n369), .A2(n368), .ZN(n448) );
  NAND2_X1 U391 ( .A1(n371), .A2(n370), .ZN(n373) );
  NAND2_X1 U392 ( .A1(n373), .A2(n372), .ZN(n447) );
  NAND2_X1 U393 ( .A1(n448), .A2(n447), .ZN(n463) );
  FA_X1 U394 ( .A(n376), .B(n375), .CI(n374), .CO(n407), .S(n385) );
  XNOR2_X1 U395 ( .A(b_in[9]), .B(a_in[5]), .ZN(n397) );
  OAI22_X1 U396 ( .A1(n487), .A2(n377), .B1(n488), .B2(n397), .ZN(n404) );
  XNOR2_X1 U397 ( .A(n378), .B(a_in[9]), .ZN(n398) );
  OAI22_X1 U398 ( .A1(n399), .A2(n379), .B1(n400), .B2(n398), .ZN(n403) );
  FA_X1 U399 ( .A(f[11]), .B(f[12]), .CI(n380), .CO(n396), .S(n374) );
  XNOR2_X1 U400 ( .A(b_in[7]), .B(a_in[7]), .ZN(n402) );
  OAI22_X1 U401 ( .A1(n420), .A2(n381), .B1(n421), .B2(n402), .ZN(n395) );
  FA_X1 U402 ( .A(n384), .B(n383), .CI(n382), .CO(n394), .S(n386) );
  FA_X1 U403 ( .A(n387), .B(n386), .CI(n385), .CO(n388), .S(n352) );
  NOR2_X1 U404 ( .A1(n389), .A2(n388), .ZN(n393) );
  INV_X1 U405 ( .A(n393), .ZN(n437) );
  NAND2_X1 U406 ( .A1(n389), .A2(n388), .ZN(n415) );
  AND2_X1 U407 ( .A1(n437), .A2(n415), .ZN(n390) );
  XNOR2_X1 U408 ( .A(n463), .B(n390), .ZN(n391) );
  AOI22_X1 U409 ( .A1(n391), .A2(n526), .B1(n509), .B2(f[13]), .ZN(n392) );
  INV_X1 U410 ( .A(n392), .ZN(n54) );
  OAI21_X1 U411 ( .B1(n463), .B2(n393), .A(n415), .ZN(n411) );
  FA_X1 U412 ( .A(n396), .B(n395), .CI(n394), .CO(n435), .S(n405) );
  XNOR2_X1 U413 ( .A(b_in[9]), .B(a_in[6]), .ZN(n416) );
  OAI22_X1 U414 ( .A1(n487), .A2(n397), .B1(n488), .B2(n416), .ZN(n426) );
  AOI21_X1 U415 ( .B1(n400), .B2(n399), .A(n398), .ZN(n401) );
  INV_X1 U416 ( .A(n401), .ZN(n429) );
  XNOR2_X1 U417 ( .A(b_in[7]), .B(a_in[8]), .ZN(n418) );
  OAI22_X1 U418 ( .A1(n420), .A2(n402), .B1(n421), .B2(n418), .ZN(n428) );
  FA_X1 U419 ( .A(n404), .B(n519), .CI(n403), .CO(n427), .S(n406) );
  FA_X1 U420 ( .A(n407), .B(n406), .CI(n405), .CO(n408), .S(n389) );
  NOR2_X1 U421 ( .A1(n409), .A2(n408), .ZN(n414) );
  INV_X1 U422 ( .A(n414), .ZN(n436) );
  NAND2_X1 U423 ( .A1(n409), .A2(n408), .ZN(n464) );
  NAND2_X1 U424 ( .A1(n436), .A2(n464), .ZN(n410) );
  XNOR2_X1 U425 ( .A(n411), .B(n410), .ZN(n412) );
  AOI22_X1 U426 ( .A1(n412), .A2(n526), .B1(n509), .B2(f[14]), .ZN(n413) );
  INV_X1 U427 ( .A(n413), .ZN(n53) );
  OR2_X1 U428 ( .A1(n415), .A2(n414), .ZN(n465) );
  XNOR2_X1 U429 ( .A(b_in[9]), .B(a_in[7]), .ZN(n423) );
  OAI22_X1 U430 ( .A1(n487), .A2(n416), .B1(n488), .B2(n423), .ZN(n425) );
  XNOR2_X1 U431 ( .A(b_in[7]), .B(a_in[9]), .ZN(n419) );
  OAI22_X1 U432 ( .A1(n420), .A2(n418), .B1(n421), .B2(n419), .ZN(n424) );
  AOI21_X1 U433 ( .B1(n421), .B2(n420), .A(n419), .ZN(n422) );
  INV_X1 U434 ( .A(n422), .ZN(n455) );
  XNOR2_X1 U435 ( .A(b_in[9]), .B(a_in[8]), .ZN(n457) );
  OAI22_X1 U436 ( .A1(n487), .A2(n423), .B1(n488), .B2(n457), .ZN(n458) );
  FA_X1 U437 ( .A(n425), .B(n518), .CI(n424), .CO(n456), .S(n432) );
  FA_X1 U438 ( .A(f[13]), .B(f[14]), .CI(n426), .CO(n431), .S(n434) );
  FA_X1 U439 ( .A(n429), .B(n428), .CI(n427), .CO(n430), .S(n433) );
  NAND2_X1 U440 ( .A1(n441), .A2(n440), .ZN(n478) );
  FA_X1 U441 ( .A(n432), .B(n431), .CI(n430), .CO(n440), .S(n439) );
  FA_X1 U442 ( .A(n435), .B(n434), .CI(n433), .CO(n438), .S(n409) );
  NAND2_X1 U443 ( .A1(n439), .A2(n438), .ZN(n472) );
  AND2_X1 U444 ( .A1(n478), .A2(n472), .ZN(n443) );
  NAND3_X1 U445 ( .A1(n465), .A2(n464), .A3(n443), .ZN(n449) );
  NAND2_X1 U446 ( .A1(n437), .A2(n436), .ZN(n462) );
  INV_X1 U447 ( .A(n462), .ZN(n445) );
  NOR2_X1 U448 ( .A1(n439), .A2(n438), .ZN(n466) );
  OR2_X1 U449 ( .A1(n441), .A2(n440), .ZN(n479) );
  INV_X1 U450 ( .A(n479), .ZN(n442) );
  AOI21_X1 U451 ( .B1(n443), .B2(n466), .A(n442), .ZN(n444) );
  OAI21_X1 U452 ( .B1(n449), .B2(n445), .A(n444), .ZN(n451) );
  INV_X1 U453 ( .A(n451), .ZN(n446) );
  NAND3_X1 U454 ( .A1(n448), .A2(n447), .A3(n446), .ZN(n453) );
  INV_X1 U455 ( .A(n449), .ZN(n450) );
  OR2_X1 U456 ( .A1(n451), .A2(n450), .ZN(n452) );
  NAND2_X1 U457 ( .A1(n453), .A2(n452), .ZN(n490) );
  FA_X1 U458 ( .A(n456), .B(n455), .CI(n454), .CO(n492), .S(n441) );
  XNOR2_X1 U459 ( .A(b_in[9]), .B(a_in[9]), .ZN(n486) );
  OAI22_X1 U460 ( .A1(n487), .A2(n457), .B1(n488), .B2(n486), .ZN(n485) );
  FA_X1 U461 ( .A(f[15]), .B(f[16]), .CI(n458), .CO(n484), .S(n454) );
  XOR2_X1 U462 ( .A(n492), .B(n491), .Z(n459) );
  XOR2_X1 U463 ( .A(n490), .B(n459), .Z(n460) );
  AOI22_X1 U464 ( .A1(n460), .A2(n526), .B1(n509), .B2(f[17]), .ZN(n461) );
  INV_X1 U465 ( .A(n461), .ZN(n50) );
  NOR2_X1 U466 ( .A1(n463), .A2(n462), .ZN(n471) );
  NAND2_X1 U467 ( .A1(n465), .A2(n464), .ZN(n475) );
  NOR2_X1 U468 ( .A1(n471), .A2(n475), .ZN(n468) );
  INV_X1 U469 ( .A(n466), .ZN(n474) );
  NAND2_X1 U470 ( .A1(n474), .A2(n472), .ZN(n467) );
  XOR2_X1 U471 ( .A(n468), .B(n467), .Z(n469) );
  AOI22_X1 U472 ( .A1(n469), .A2(n526), .B1(n509), .B2(f[15]), .ZN(n470) );
  INV_X1 U473 ( .A(n470), .ZN(n52) );
  NAND2_X1 U474 ( .A1(n471), .A2(n474), .ZN(n477) );
  INV_X1 U475 ( .A(n472), .ZN(n473) );
  AOI21_X1 U476 ( .B1(n475), .B2(n474), .A(n473), .ZN(n476) );
  NAND2_X1 U477 ( .A1(n477), .A2(n476), .ZN(n481) );
  NAND2_X1 U478 ( .A1(n479), .A2(n478), .ZN(n480) );
  XNOR2_X1 U479 ( .A(n481), .B(n480), .ZN(n482) );
  AOI22_X1 U480 ( .A1(n482), .A2(n526), .B1(n509), .B2(f[16]), .ZN(n483) );
  INV_X1 U481 ( .A(n483), .ZN(n51) );
  FA_X1 U482 ( .A(n485), .B(n517), .CI(n484), .CO(n508), .S(n491) );
  AOI21_X1 U483 ( .B1(n488), .B2(n487), .A(n486), .ZN(n489) );
  INV_X1 U484 ( .A(n489), .ZN(n496) );
  NAND2_X1 U485 ( .A1(n490), .A2(n492), .ZN(n495) );
  NAND2_X1 U486 ( .A1(n490), .A2(n491), .ZN(n494) );
  NAND2_X1 U487 ( .A1(n492), .A2(n491), .ZN(n493) );
  NAND3_X1 U488 ( .A1(n495), .A2(n494), .A3(n493), .ZN(n506) );
  FA_X1 U489 ( .A(f[17]), .B(f[18]), .CI(n496), .CO(n497), .S(n507) );
  XNOR2_X1 U490 ( .A(n516), .B(n497), .ZN(n498) );
  XNOR2_X1 U491 ( .A(n499), .B(n498), .ZN(n500) );
  NAND2_X1 U492 ( .A1(n500), .A2(n526), .ZN(n502) );
  NAND2_X1 U493 ( .A1(n509), .A2(f[19]), .ZN(n501) );
  NAND2_X1 U494 ( .A1(n502), .A2(n501), .ZN(n48) );
  AOI22_X1 U495 ( .A1(n514), .A2(b[9]), .B1(n513), .B2(b_in[9]), .ZN(n503) );
  INV_X1 U496 ( .A(n503), .ZN(n68) );
  AOI22_X1 U497 ( .A1(n514), .A2(b[1]), .B1(n513), .B2(b_in[1]), .ZN(n504) );
  INV_X1 U498 ( .A(n504), .ZN(n76) );
  AOI22_X1 U499 ( .A1(n514), .A2(b[7]), .B1(n513), .B2(b_in[7]), .ZN(n505) );
  INV_X1 U500 ( .A(n505), .ZN(n70) );
  FA_X1 U501 ( .A(n508), .B(n507), .CI(n506), .CO(n499), .S(n510) );
  AOI22_X1 U502 ( .A1(n510), .A2(n526), .B1(n509), .B2(f[18]), .ZN(n511) );
  INV_X1 U503 ( .A(n511), .ZN(n49) );
  AOI22_X1 U504 ( .A1(n514), .A2(b[3]), .B1(n513), .B2(b_in[3]), .ZN(n512) );
  INV_X1 U505 ( .A(n512), .ZN(n74) );
  AOI22_X1 U506 ( .A1(n514), .A2(b[5]), .B1(n513), .B2(b_in[5]), .ZN(n515) );
  INV_X1 U507 ( .A(n515), .ZN(n72) );
endmodule

