
module part2_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   N46, N47, N55, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n101, n102, n105, n106,
         n109, n112, n113, n115, n116, n117, \DP_OP_37J1_122_8065/n409 , n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796;
  wire   [9:0] a_in;
  wire   [9:0] b_in;
  assign f[19] = N55;

  DFF_X1 enable_f_reg ( .D(n796), .CK(clk), .QN(n768) );
  DFF_X1 valid_out_reg ( .D(n795), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[19]  ( .D(n78), .CK(clk), .Q(N55), .QN(n769) );
  DFF_X1 \f_reg[17]  ( .D(n80), .CK(clk), .Q(f[17]), .QN(n773) );
  DFF_X1 \f_reg[10]  ( .D(n87), .CK(clk), .Q(f[10]), .QN(n774) );
  DFF_X1 \f_reg[1]  ( .D(n96), .CK(clk), .Q(f[1]), .QN(n783) );
  DFF_X1 \a_in_reg[8]  ( .D(n116), .CK(clk), .Q(a_in[8]), .QN(n750) );
  DFF_X1 \a_in_reg[7]  ( .D(n115), .CK(clk), .Q(a_in[7]), .QN(n753) );
  DFF_X1 \a_in_reg[5]  ( .D(n113), .CK(clk), .Q(a_in[5]) );
  DFF_X1 \a_in_reg[4]  ( .D(n112), .CK(clk), .Q(a_in[4]), .QN(n751) );
  DFF_X1 \b_in_reg[8]  ( .D(n106), .CK(clk), .Q(b_in[8]), .QN(n755) );
  DFF_X1 \b_in_reg[4]  ( .D(n102), .CK(clk), .Q(b_in[4]), .QN(n758) );
  DFF_X1 \b_in_reg[7]  ( .D(n105), .CK(clk), .Q(b_in[7]), .QN(n754) );
  DFF_X1 \b_in_reg[3]  ( .D(n101), .CK(clk), .Q(b_in[3]), .QN(n759) );
  DFF_X1 \b_in_reg[1]  ( .D(n786), .CK(clk), .Q(n757), .QN(
        \DP_OP_37J1_122_8065/n409 ) );
  DFF_X1 \b_in_reg[5]  ( .D(n785), .CK(clk), .Q(n756), .QN(b_in[5]) );
  DFF_X1 \b_in_reg[9]  ( .D(n791), .CK(clk), .Q(n766), .QN(N47) );
  DFF_X1 \b_in_reg[6]  ( .D(n792), .CK(clk), .Q(n761), .QN(b_in[6]) );
  DFF_X1 \b_in_reg[2]  ( .D(n793), .CK(clk), .Q(n760), .QN(b_in[2]) );
  DFF_X1 \a_in_reg[9]  ( .D(n117), .CK(clk), .Q(N46), .QN(n752) );
  DFF_X2 \f_reg[5]  ( .D(n92), .CK(clk), .Q(f[5]), .QN(n776) );
  DFF_X2 \f_reg[6]  ( .D(n91), .CK(clk), .Q(f[6]), .QN(n780) );
  DFF_X2 \f_reg[18]  ( .D(n79), .CK(clk), .Q(f[18]), .QN(n784) );
  DFF_X2 \f_reg[7]  ( .D(n90), .CK(clk), .Q(f[7]), .QN(n763) );
  DFF_X2 \f_reg[9]  ( .D(n88), .CK(clk), .Q(f[9]), .QN(n762) );
  DFF_X2 \f_reg[13]  ( .D(n84), .CK(clk), .Q(f[13]), .QN(n764) );
  DFF_X1 \a_in_reg[2]  ( .D(n789), .CK(clk), .QN(a_in[2]) );
  DFF_X1 \a_in_reg[3]  ( .D(n788), .CK(clk), .QN(a_in[3]) );
  DFF_X1 \a_in_reg[0]  ( .D(n790), .CK(clk), .QN(a_in[0]) );
  DFF_X1 \b_in_reg[0]  ( .D(n794), .CK(clk), .Q(n765), .QN(b_in[0]) );
  DFF_X1 \a_in_reg[6]  ( .D(n787), .CK(clk), .QN(a_in[6]) );
  DFF_X2 \f_reg[0]  ( .D(n97), .CK(clk), .Q(f[0]), .QN(n767) );
  DFF_X2 \f_reg[3]  ( .D(n94), .CK(clk), .Q(f[3]), .QN(n775) );
  DFF_X2 \f_reg[4]  ( .D(n93), .CK(clk), .Q(f[4]), .QN(n779) );
  DFF_X2 \f_reg[8]  ( .D(n89), .CK(clk), .Q(f[8]), .QN(n778) );
  DFF_X2 \f_reg[11]  ( .D(n86), .CK(clk), .Q(f[11]), .QN(n771) );
  DFF_X2 \f_reg[16]  ( .D(n81), .CK(clk), .Q(f[16]), .QN(n781) );
  DFF_X2 \f_reg[2]  ( .D(n95), .CK(clk), .Q(f[2]), .QN(n770) );
  DFF_X2 \f_reg[14]  ( .D(n83), .CK(clk), .Q(f[14]), .QN(n777) );
  DFF_X2 \f_reg[15]  ( .D(n82), .CK(clk), .Q(f[15]), .QN(n772) );
  DFF_X1 \a_in_reg[1]  ( .D(n109), .CK(clk), .Q(a_in[1]), .QN(n140) );
  DFF_X1 \f_reg[12]  ( .D(n85), .CK(clk), .Q(f[12]), .QN(n782) );
  NAND3_X1 U122 ( .A1(n229), .A2(n230), .A3(n228), .ZN(n426) );
  XNOR2_X2 U123 ( .A(n214), .B(n265), .ZN(n270) );
  XNOR2_X1 U124 ( .A(n118), .B(n164), .ZN(n735) );
  AOI21_X1 U125 ( .B1(n617), .B2(n618), .A(n616), .ZN(n118) );
  NOR2_X1 U126 ( .A1(n119), .A2(n728), .ZN(n612) );
  NAND2_X1 U127 ( .A1(n121), .A2(n120), .ZN(n119) );
  NOR2_X1 U128 ( .A1(n727), .A2(n495), .ZN(n120) );
  INV_X1 U129 ( .A(n726), .ZN(n121) );
  BUF_X1 U130 ( .A(\DP_OP_37J1_122_8065/n409 ), .Z(n628) );
  BUF_X2 U131 ( .A(b_in[7]), .Z(n746) );
  AND3_X2 U132 ( .A1(n139), .A2(n732), .A3(n731), .ZN(n611) );
  CLKBUF_X1 U133 ( .A(n535), .Z(n158) );
  AND2_X1 U134 ( .A1(n713), .A2(n144), .ZN(n697) );
  BUF_X1 U135 ( .A(n731), .Z(n667) );
  AOI21_X1 U136 ( .B1(n497), .B2(n544), .A(n496), .ZN(n498) );
  OR2_X1 U137 ( .A1(n479), .A2(n480), .ZN(n544) );
  OR2_X1 U138 ( .A1(n385), .A2(n384), .ZN(n558) );
  NAND2_X1 U139 ( .A1(n123), .A2(n122), .ZN(n384) );
  NAND2_X1 U140 ( .A1(n357), .A2(n124), .ZN(n123) );
  NAND2_X1 U141 ( .A1(n126), .A2(n125), .ZN(n124) );
  OAI21_X1 U142 ( .B1(n570), .B2(n573), .A(n571), .ZN(n577) );
  INV_X1 U143 ( .A(n359), .ZN(n126) );
  NAND2_X1 U144 ( .A1(n359), .A2(n358), .ZN(n122) );
  INV_X1 U145 ( .A(n358), .ZN(n125) );
  NAND2_X1 U146 ( .A1(n130), .A2(n129), .ZN(n232) );
  OAI21_X1 U147 ( .B1(n242), .B2(f[8]), .A(n131), .ZN(n130) );
  OR2_X1 U148 ( .A1(n213), .A2(f[10]), .ZN(n284) );
  BUF_X1 U149 ( .A(n436), .Z(n153) );
  INV_X1 U150 ( .A(n141), .ZN(n526) );
  INV_X1 U151 ( .A(n750), .ZN(n722) );
  XOR2_X1 U152 ( .A(n759), .B(a_in[8]), .Z(n206) );
  XNOR2_X1 U153 ( .A(n213), .B(f[10]), .ZN(n226) );
  OAI22_X1 U154 ( .A1(n437), .A2(n203), .B1(n204), .B2(n436), .ZN(n213) );
  BUF_X2 U155 ( .A(n205), .Z(n244) );
  XNOR2_X1 U156 ( .A(n357), .B(n127), .ZN(n342) );
  XNOR2_X1 U157 ( .A(n359), .B(n358), .ZN(n127) );
  NAND2_X1 U158 ( .A1(n535), .A2(n432), .ZN(n434) );
  NOR2_X1 U159 ( .A1(n253), .A2(n594), .ZN(n535) );
  XNOR2_X1 U160 ( .A(n128), .B(n131), .ZN(n405) );
  OAI22_X1 U161 ( .A1(n371), .A2(n369), .B1(n222), .B2(n765), .ZN(n131) );
  XNOR2_X1 U162 ( .A(n242), .B(f[8]), .ZN(n128) );
  NAND2_X1 U163 ( .A1(n242), .A2(f[8]), .ZN(n129) );
  XNOR2_X1 U164 ( .A(n531), .B(n132), .ZN(n139) );
  INV_X1 U165 ( .A(n530), .ZN(n132) );
  NAND2_X1 U166 ( .A1(n617), .A2(n614), .ZN(n531) );
  NAND2_X1 U167 ( .A1(n138), .A2(n133), .ZN(n617) );
  AND2_X1 U168 ( .A1(n517), .A2(n521), .ZN(n133) );
  OAI21_X1 U169 ( .B1(n504), .B2(n434), .A(n433), .ZN(n138) );
  BUF_X1 U170 ( .A(n728), .Z(n134) );
  XNOR2_X1 U171 ( .A(n272), .B(n271), .ZN(n135) );
  XNOR2_X1 U172 ( .A(n135), .B(n270), .ZN(n136) );
  AOI21_X1 U173 ( .B1(n546), .B2(n423), .A(n422), .ZN(n137) );
  XNOR2_X1 U174 ( .A(n757), .B(n140), .ZN(n313) );
  XOR2_X1 U175 ( .A(n754), .B(n755), .Z(n141) );
  BUF_X1 U176 ( .A(n726), .Z(n142) );
  BUF_X1 U177 ( .A(n191), .Z(n143) );
  OR2_X1 U178 ( .A1(n740), .A2(n776), .ZN(n144) );
  AND2_X1 U179 ( .A1(n713), .A2(n145), .ZN(n700) );
  OR2_X1 U180 ( .A1(n740), .A2(n763), .ZN(n145) );
  AND2_X1 U181 ( .A1(n713), .A2(n146), .ZN(n694) );
  OR2_X1 U182 ( .A1(n740), .A2(n780), .ZN(n146) );
  AND2_X1 U183 ( .A1(n713), .A2(n181), .ZN(n703) );
  NAND2_X1 U184 ( .A1(n660), .A2(n659), .ZN(n147) );
  NAND2_X1 U185 ( .A1(n660), .A2(n659), .ZN(n148) );
  NAND2_X1 U186 ( .A1(n660), .A2(n659), .ZN(n709) );
  BUF_X1 U187 ( .A(n289), .Z(n149) );
  NAND2_X1 U188 ( .A1(n195), .A2(n186), .ZN(n150) );
  OAI22_X1 U189 ( .A1(n150), .A2(n211), .B1(n526), .B2(n261), .ZN(n151) );
  XNOR2_X1 U190 ( .A(n754), .B(n755), .ZN(n195) );
  NOR2_X1 U191 ( .A1(n511), .A2(n510), .ZN(n152) );
  XOR2_X1 U192 ( .A(n757), .B(a_in[8]), .Z(n222) );
  NAND2_X1 U193 ( .A1(n185), .A2(n184), .ZN(n154) );
  NAND2_X1 U194 ( .A1(n185), .A2(n184), .ZN(n155) );
  BUF_X1 U195 ( .A(n134), .Z(n156) );
  NAND2_X1 U196 ( .A1(n185), .A2(n184), .ZN(n470) );
  OAI211_X1 U197 ( .C1(n388), .C2(n387), .A(n589), .B(n386), .ZN(n157) );
  NAND2_X1 U198 ( .A1(n274), .A2(n273), .ZN(n428) );
  NAND2_X1 U199 ( .A1(n278), .A2(n277), .ZN(n445) );
  NAND2_X1 U200 ( .A1(f[11]), .A2(f[12]), .ZN(n277) );
  NAND2_X1 U201 ( .A1(n276), .A2(n275), .ZN(n278) );
  NAND2_X1 U202 ( .A1(n771), .A2(n782), .ZN(n275) );
  INV_X1 U203 ( .A(n537), .ZN(n506) );
  NAND2_X1 U204 ( .A1(n394), .A2(n393), .ZN(n395) );
  INV_X1 U205 ( .A(n397), .ZN(n393) );
  NAND2_X1 U206 ( .A1(n417), .A2(n416), .ZN(n418) );
  NAND2_X1 U207 ( .A1(n410), .A2(n415), .ZN(n416) );
  NAND2_X1 U208 ( .A1(n414), .A2(n413), .ZN(n417) );
  NAND2_X1 U209 ( .A1(n412), .A2(n411), .ZN(n413) );
  AND2_X1 U210 ( .A1(n366), .A2(f[7]), .ZN(n406) );
  INV_X1 U211 ( .A(n460), .ZN(n456) );
  XNOR2_X1 U212 ( .A(n445), .B(n444), .ZN(n283) );
  NAND2_X1 U213 ( .A1(n267), .A2(n266), .ZN(n268) );
  CLKBUF_X1 U214 ( .A(n505), .Z(n536) );
  INV_X1 U215 ( .A(n410), .ZN(n412) );
  INV_X1 U216 ( .A(n415), .ZN(n411) );
  XNOR2_X1 U217 ( .A(n276), .B(n256), .ZN(n287) );
  XNOR2_X1 U218 ( .A(f[11]), .B(f[12]), .ZN(n256) );
  AND2_X1 U219 ( .A1(n305), .A2(f[3]), .ZN(n338) );
  NAND2_X1 U220 ( .A1(n400), .A2(n399), .ZN(n409) );
  NAND2_X1 U221 ( .A1(n396), .A2(n395), .ZN(n400) );
  NAND2_X1 U222 ( .A1(n378), .A2(n377), .ZN(n382) );
  NAND2_X1 U223 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U224 ( .A1(n374), .A2(n373), .ZN(n378) );
  OR2_X1 U225 ( .A1(n376), .A2(n375), .ZN(n373) );
  XNOR2_X1 U226 ( .A(n396), .B(n372), .ZN(n414) );
  XNOR2_X1 U227 ( .A(n374), .B(n356), .ZN(n385) );
  XNOR2_X1 U228 ( .A(n376), .B(n375), .ZN(n356) );
  NAND2_X1 U229 ( .A1(n340), .A2(n339), .ZN(n341) );
  NAND2_X1 U230 ( .A1(n338), .A2(n337), .ZN(n339) );
  NAND2_X1 U231 ( .A1(n336), .A2(n335), .ZN(n340) );
  OR2_X1 U232 ( .A1(n338), .A2(n337), .ZN(n335) );
  XNOR2_X1 U233 ( .A(n336), .B(n300), .ZN(n325) );
  XNOR2_X1 U234 ( .A(n338), .B(n337), .ZN(n300) );
  NAND2_X1 U235 ( .A1(n391), .A2(n165), .ZN(n248) );
  NAND2_X1 U236 ( .A1(n463), .A2(n462), .ZN(n477) );
  NAND2_X1 U237 ( .A1(n461), .A2(n460), .ZN(n462) );
  NAND2_X1 U238 ( .A1(n459), .A2(n458), .ZN(n463) );
  NAND2_X1 U239 ( .A1(n445), .A2(n444), .ZN(n447) );
  BUF_X1 U240 ( .A(n547), .Z(n548) );
  BUF_X1 U241 ( .A(n549), .Z(n602) );
  CLKBUF_X1 U242 ( .A(n596), .Z(n597) );
  INV_X1 U243 ( .A(n540), .ZN(n497) );
  XNOR2_X1 U244 ( .A(n515), .B(n514), .ZN(n727) );
  OAI21_X1 U245 ( .B1(n504), .B2(n509), .A(n508), .ZN(n515) );
  XNOR2_X1 U246 ( .A(n538), .B(n163), .ZN(n708) );
  BUF_X1 U247 ( .A(n533), .Z(n534) );
  BUF_X1 U248 ( .A(n629), .Z(n743) );
  NAND2_X1 U249 ( .A1(n768), .A2(n716), .ZN(n740) );
  NOR2_X1 U250 ( .A1(n768), .A2(reset), .ZN(n795) );
  AND2_X1 U251 ( .A1(valid_in), .A2(n716), .ZN(n796) );
  AND2_X1 U252 ( .A1(n210), .A2(f[9]), .ZN(n159) );
  BUF_X1 U253 ( .A(b_in[5]), .Z(n329) );
  XOR2_X1 U254 ( .A(n746), .B(a_in[0]), .Z(n160) );
  AND2_X1 U255 ( .A1(n521), .A2(n519), .ZN(n161) );
  AND2_X1 U256 ( .A1(n544), .A2(n543), .ZN(n162) );
  AND2_X1 U257 ( .A1(n507), .A2(n537), .ZN(n163) );
  NAND2_X1 U258 ( .A1(n622), .A2(n621), .ZN(n164) );
  OR2_X1 U259 ( .A1(n389), .A2(n390), .ZN(n165) );
  OR2_X1 U260 ( .A1(n740), .A2(n770), .ZN(n166) );
  OR2_X1 U261 ( .A1(n740), .A2(n767), .ZN(n167) );
  OR2_X1 U262 ( .A1(n740), .A2(n775), .ZN(n168) );
  OR2_X1 U263 ( .A1(n740), .A2(n772), .ZN(n169) );
  OR2_X1 U264 ( .A1(n740), .A2(n783), .ZN(n170) );
  OR2_X1 U265 ( .A1(n740), .A2(n779), .ZN(n171) );
  OR2_X1 U266 ( .A1(n740), .A2(n774), .ZN(n172) );
  OR2_X1 U267 ( .A1(n740), .A2(n777), .ZN(n173) );
  OR2_X1 U268 ( .A1(n740), .A2(n778), .ZN(n174) );
  OR2_X1 U269 ( .A1(n740), .A2(n771), .ZN(n175) );
  OR2_X1 U270 ( .A1(n740), .A2(n773), .ZN(n176) );
  OR2_X1 U271 ( .A1(n740), .A2(n781), .ZN(n177) );
  OR2_X1 U272 ( .A1(n740), .A2(n762), .ZN(n178) );
  OR2_X1 U273 ( .A1(n740), .A2(n782), .ZN(n179) );
  OR2_X1 U274 ( .A1(n740), .A2(n764), .ZN(n180) );
  OR2_X1 U275 ( .A1(n740), .A2(n784), .ZN(n181) );
  OR2_X2 U276 ( .A1(n757), .A2(b_in[0]), .ZN(n371) );
  XNOR2_X1 U277 ( .A(n757), .B(n752), .ZN(n188) );
  AOI21_X1 U278 ( .B1(n371), .B2(n765), .A(n188), .ZN(n182) );
  INV_X1 U279 ( .A(n182), .ZN(n209) );
  XNOR2_X1 U280 ( .A(b_in[3]), .B(n760), .ZN(n183) );
  XNOR2_X1 U281 ( .A(b_in[2]), .B(\DP_OP_37J1_122_8065/n409 ), .ZN(n191) );
  NAND2_X1 U282 ( .A1(n183), .A2(n191), .ZN(n205) );
  BUF_X4 U283 ( .A(b_in[3]), .Z(n629) );
  XNOR2_X1 U284 ( .A(n629), .B(a_in[7]), .ZN(n192) );
  OAI22_X1 U285 ( .A1(n192), .A2(n205), .B1(n143), .B2(n206), .ZN(n208) );
  XNOR2_X1 U286 ( .A(b_in[5]), .B(b_in[6]), .ZN(n185) );
  XNOR2_X1 U287 ( .A(b_in[7]), .B(n761), .ZN(n184) );
  XNOR2_X1 U288 ( .A(n746), .B(a_in[3]), .ZN(n193) );
  XNOR2_X1 U289 ( .A(b_in[5]), .B(b_in[6]), .ZN(n353) );
  BUF_X2 U290 ( .A(n353), .Z(n471) );
  XNOR2_X1 U291 ( .A(n754), .B(n751), .ZN(n202) );
  OAI22_X1 U292 ( .A1(n470), .A2(n193), .B1(n471), .B2(n202), .ZN(n207) );
  XOR2_X1 U293 ( .A(b_in[8]), .B(N47), .Z(n186) );
  NAND2_X1 U294 ( .A1(n186), .A2(n195), .ZN(n201) );
  OR2_X1 U295 ( .A1(a_in[0]), .A2(n766), .ZN(n187) );
  OAI22_X1 U296 ( .A1(n201), .A2(n766), .B1(n187), .B2(n195), .ZN(n225) );
  BUF_X2 U297 ( .A(\DP_OP_37J1_122_8065/n409 ), .Z(n748) );
  OAI22_X1 U298 ( .A1(n371), .A2(n222), .B1(n188), .B2(n765), .ZN(n224) );
  XNOR2_X1 U299 ( .A(n759), .B(n758), .ZN(n190) );
  XNOR2_X1 U300 ( .A(b_in[4]), .B(n756), .ZN(n189) );
  NAND2_X2 U301 ( .A1(n189), .A2(n190), .ZN(n437) );
  BUF_X2 U302 ( .A(b_in[5]), .Z(n745) );
  XNOR2_X1 U303 ( .A(n745), .B(a_in[4]), .ZN(n221) );
  BUF_X2 U304 ( .A(n190), .Z(n436) );
  XNOR2_X1 U305 ( .A(n329), .B(a_in[5]), .ZN(n203) );
  OAI22_X1 U306 ( .A1(n437), .A2(n221), .B1(n436), .B2(n203), .ZN(n223) );
  BUF_X2 U307 ( .A(n205), .Z(n348) );
  XNOR2_X1 U308 ( .A(n629), .B(a_in[6]), .ZN(n220) );
  INV_X1 U309 ( .A(n191), .ZN(n309) );
  OAI22_X1 U310 ( .A1(n348), .A2(n220), .B1(n143), .B2(n192), .ZN(n234) );
  XNOR2_X1 U311 ( .A(n746), .B(a_in[2]), .ZN(n219) );
  OAI22_X1 U312 ( .A1(n471), .A2(n193), .B1(n155), .B2(n219), .ZN(n235) );
  OR2_X1 U313 ( .A1(n234), .A2(n235), .ZN(n198) );
  INV_X1 U314 ( .A(N47), .ZN(n194) );
  INV_X2 U315 ( .A(n194), .ZN(n486) );
  XNOR2_X1 U316 ( .A(n486), .B(a_in[0]), .ZN(n197) );
  XOR2_X1 U317 ( .A(n766), .B(a_in[1]), .Z(n212) );
  OR2_X1 U318 ( .A1(n212), .A2(n195), .ZN(n196) );
  OAI21_X1 U319 ( .B1(n201), .B2(n197), .A(n196), .ZN(n210) );
  XNOR2_X1 U320 ( .A(n210), .B(n762), .ZN(n237) );
  NAND2_X1 U321 ( .A1(n198), .A2(n237), .ZN(n200) );
  NAND2_X1 U322 ( .A1(n235), .A2(n234), .ZN(n199) );
  NAND2_X1 U323 ( .A1(n200), .A2(n199), .ZN(n216) );
  XNOR2_X1 U324 ( .A(n486), .B(a_in[2]), .ZN(n211) );
  XNOR2_X1 U325 ( .A(n486), .B(a_in[3]), .ZN(n261) );
  OAI22_X1 U326 ( .A1(n150), .A2(n211), .B1(n526), .B2(n261), .ZN(n286) );
  XNOR2_X1 U327 ( .A(n746), .B(a_in[5]), .ZN(n262) );
  OAI22_X1 U328 ( .A1(n471), .A2(n262), .B1(n155), .B2(n202), .ZN(n285) );
  XNOR2_X1 U329 ( .A(n329), .B(a_in[6]), .ZN(n204) );
  XNOR2_X1 U330 ( .A(n272), .B(n271), .ZN(n215) );
  XNOR2_X1 U331 ( .A(n756), .B(n753), .ZN(n255) );
  OAI22_X1 U332 ( .A1(n437), .A2(n204), .B1(n436), .B2(n255), .ZN(n258) );
  XNOR2_X1 U333 ( .A(n629), .B(N46), .ZN(n263) );
  OAI22_X1 U334 ( .A1(n244), .A2(n206), .B1(n333), .B2(n263), .ZN(n257) );
  FA_X1 U335 ( .A(n209), .B(n208), .CI(n207), .CO(n266), .S(n218) );
  XNOR2_X1 U336 ( .A(n267), .B(n266), .ZN(n214) );
  OAI22_X1 U337 ( .A1(n150), .A2(n212), .B1(n526), .B2(n211), .ZN(n227) );
  XNOR2_X1 U338 ( .A(n215), .B(n270), .ZN(n427) );
  FA_X1 U339 ( .A(n218), .B(n217), .CI(n216), .CO(n272), .S(n251) );
  XNOR2_X1 U340 ( .A(n746), .B(a_in[1]), .ZN(n239) );
  OAI22_X1 U341 ( .A1(n154), .A2(n239), .B1(n471), .B2(n219), .ZN(n403) );
  XNOR2_X1 U342 ( .A(n629), .B(a_in[5]), .ZN(n243) );
  INV_X1 U343 ( .A(n309), .ZN(n346) );
  OAI22_X1 U344 ( .A1(n244), .A2(n243), .B1(n346), .B2(n220), .ZN(n402) );
  XNOR2_X1 U345 ( .A(n745), .B(a_in[3]), .ZN(n245) );
  OAI22_X1 U346 ( .A1(n437), .A2(n245), .B1(n436), .B2(n221), .ZN(n401) );
  AND2_X1 U347 ( .A1(a_in[0]), .A2(n141), .ZN(n242) );
  XNOR2_X1 U348 ( .A(n628), .B(a_in[7]), .ZN(n369) );
  FA_X1 U349 ( .A(n225), .B(n224), .CI(n223), .CO(n217), .S(n231) );
  NAND2_X1 U350 ( .A1(n251), .A2(n250), .ZN(n230) );
  FA_X1 U351 ( .A(n159), .B(n227), .CI(n226), .CO(n265), .S(n249) );
  NAND2_X1 U352 ( .A1(n251), .A2(n249), .ZN(n229) );
  NAND2_X1 U353 ( .A1(n250), .A2(n249), .ZN(n228) );
  NOR2_X1 U354 ( .A1(n136), .A2(n426), .ZN(n253) );
  FA_X1 U355 ( .A(n233), .B(n232), .CI(n231), .CO(n250), .S(n391) );
  XNOR2_X1 U356 ( .A(n234), .B(n235), .ZN(n236) );
  XNOR2_X1 U357 ( .A(n237), .B(n236), .ZN(n389) );
  INV_X1 U358 ( .A(n155), .ZN(n238) );
  NAND2_X1 U359 ( .A1(n238), .A2(n160), .ZN(n241) );
  OR2_X1 U360 ( .A1(n471), .A2(n239), .ZN(n240) );
  NAND2_X1 U361 ( .A1(n241), .A2(n240), .ZN(n366) );
  XNOR2_X1 U362 ( .A(n629), .B(a_in[4]), .ZN(n345) );
  INV_X1 U363 ( .A(n309), .ZN(n333) );
  OAI22_X1 U364 ( .A1(n244), .A2(n345), .B1(n333), .B2(n243), .ZN(n365) );
  XNOR2_X1 U365 ( .A(n745), .B(a_in[2]), .ZN(n343) );
  OAI22_X1 U366 ( .A1(n437), .A2(n343), .B1(n436), .B2(n245), .ZN(n364) );
  OR2_X1 U367 ( .A1(a_in[0]), .A2(n754), .ZN(n246) );
  OAI22_X1 U368 ( .A1(n246), .A2(n471), .B1(n154), .B2(n754), .ZN(n363) );
  NAND2_X1 U369 ( .A1(n390), .A2(n389), .ZN(n247) );
  NAND2_X1 U370 ( .A1(n248), .A2(n247), .ZN(n424) );
  XNOR2_X1 U371 ( .A(n250), .B(n249), .ZN(n252) );
  XNOR2_X1 U372 ( .A(n252), .B(n251), .ZN(n425) );
  NOR2_X1 U373 ( .A1(n424), .A2(n425), .ZN(n594) );
  XNOR2_X1 U374 ( .A(n329), .B(n722), .ZN(n291) );
  OR2_X1 U375 ( .A1(n291), .A2(n436), .ZN(n254) );
  OAI21_X1 U376 ( .B1(n437), .B2(n255), .A(n254), .ZN(n276) );
  FA_X1 U377 ( .A(n258), .B(n771), .CI(n257), .CO(n289), .S(n267) );
  XNOR2_X1 U378 ( .A(n289), .B(n287), .ZN(n259) );
  FA_X1 U379 ( .A(n151), .B(n285), .CI(n284), .CO(n290) );
  XNOR2_X1 U380 ( .A(n259), .B(n290), .ZN(n297) );
  XNOR2_X1 U381 ( .A(n486), .B(a_in[4]), .ZN(n279) );
  OR2_X1 U382 ( .A1(n526), .A2(n279), .ZN(n260) );
  OAI21_X1 U383 ( .B1(n150), .B2(n261), .A(n260), .ZN(n282) );
  XNOR2_X1 U384 ( .A(n746), .B(a_in[6]), .ZN(n292) );
  OAI22_X1 U385 ( .A1(n154), .A2(n262), .B1(n471), .B2(n292), .ZN(n281) );
  AOI21_X1 U386 ( .B1(n346), .B2(n348), .A(n263), .ZN(n264) );
  INV_X1 U387 ( .A(n264), .ZN(n280) );
  OAI21_X1 U388 ( .B1(n267), .B2(n266), .A(n265), .ZN(n269) );
  NAND2_X1 U389 ( .A1(n269), .A2(n268), .ZN(n295) );
  OAI21_X1 U390 ( .B1(n272), .B2(n271), .A(n270), .ZN(n274) );
  NAND2_X1 U391 ( .A1(n272), .A2(n271), .ZN(n273) );
  NOR2_X1 U392 ( .A1(n429), .A2(n428), .ZN(n505) );
  XNOR2_X1 U393 ( .A(n486), .B(a_in[5]), .ZN(n439) );
  OAI22_X1 U394 ( .A1(n150), .A2(n279), .B1(n526), .B2(n439), .ZN(n444) );
  FA_X1 U395 ( .A(n282), .B(n281), .CI(n280), .CO(n443), .S(n296) );
  XNOR2_X1 U396 ( .A(n283), .B(n443), .ZN(n459) );
  FA_X1 U397 ( .A(n286), .B(n285), .CI(n284), .CO(n288), .S(n271) );
  OAI21_X1 U398 ( .B1(n288), .B2(n149), .A(n287), .ZN(n455) );
  NAND2_X1 U399 ( .A1(n290), .A2(n149), .ZN(n454) );
  NAND2_X1 U400 ( .A1(n455), .A2(n454), .ZN(n293) );
  XNOR2_X1 U401 ( .A(n745), .B(N46), .ZN(n435) );
  OAI22_X1 U402 ( .A1(n437), .A2(n291), .B1(n436), .B2(n435), .ZN(n441) );
  XNOR2_X1 U403 ( .A(n746), .B(a_in[7]), .ZN(n442) );
  OAI22_X1 U404 ( .A1(n471), .A2(n442), .B1(n154), .B2(n292), .ZN(n440) );
  XNOR2_X1 U405 ( .A(n293), .B(n460), .ZN(n294) );
  XNOR2_X1 U406 ( .A(n294), .B(n459), .ZN(n511) );
  FA_X1 U407 ( .A(n297), .B(n296), .CI(n295), .CO(n510), .S(n429) );
  NOR2_X1 U408 ( .A1(n511), .A2(n510), .ZN(n430) );
  NOR2_X1 U409 ( .A1(n505), .A2(n430), .ZN(n432) );
  INV_X1 U410 ( .A(n436), .ZN(n298) );
  AND2_X1 U411 ( .A1(a_in[0]), .A2(n298), .ZN(n327) );
  XNOR2_X1 U412 ( .A(n748), .B(a_in[3]), .ZN(n299) );
  XNOR2_X1 U413 ( .A(n748), .B(a_in[4]), .ZN(n332) );
  OAI22_X1 U414 ( .A1(n371), .A2(n299), .B1(n332), .B2(n765), .ZN(n326) );
  XNOR2_X1 U415 ( .A(n628), .B(a_in[2]), .ZN(n310) );
  OAI22_X1 U416 ( .A1(n310), .A2(n371), .B1(n299), .B2(n765), .ZN(n305) );
  XNOR2_X1 U417 ( .A(n629), .B(a_in[1]), .ZN(n303) );
  XNOR2_X1 U418 ( .A(n629), .B(a_in[2]), .ZN(n334) );
  OAI22_X1 U419 ( .A1(n348), .A2(n303), .B1(n346), .B2(n334), .ZN(n337) );
  INV_X1 U420 ( .A(n629), .ZN(n302) );
  OR2_X1 U421 ( .A1(a_in[0]), .A2(n302), .ZN(n301) );
  OAI22_X1 U422 ( .A1(n348), .A2(n302), .B1(n301), .B2(n346), .ZN(n308) );
  XNOR2_X1 U423 ( .A(n629), .B(a_in[0]), .ZN(n304) );
  OAI22_X1 U424 ( .A1(n348), .A2(n304), .B1(n333), .B2(n303), .ZN(n307) );
  XNOR2_X1 U425 ( .A(n305), .B(n775), .ZN(n306) );
  NOR2_X1 U426 ( .A1(n325), .A2(n324), .ZN(n565) );
  FA_X1 U427 ( .A(n308), .B(n307), .CI(n306), .CO(n324), .S(n322) );
  AND2_X1 U428 ( .A1(n309), .A2(a_in[0]), .ZN(n312) );
  OAI22_X1 U429 ( .A1(n371), .A2(n313), .B1(n310), .B2(n765), .ZN(n311) );
  OR2_X1 U430 ( .A1(n322), .A2(n321), .ZN(n576) );
  FA_X1 U431 ( .A(n312), .B(f[2]), .CI(n311), .CO(n321), .S(n320) );
  OAI22_X1 U432 ( .A1(n371), .A2(a_in[0]), .B1(n313), .B2(n765), .ZN(n314) );
  NOR2_X1 U433 ( .A1(n320), .A2(n319), .ZN(n570) );
  HA_X1 U434 ( .A(n314), .B(f[1]), .CO(n319), .S(n317) );
  OR2_X1 U435 ( .A1(a_in[0]), .A2(n757), .ZN(n315) );
  NAND2_X1 U436 ( .A1(n315), .A2(n371), .ZN(n316) );
  NOR2_X1 U437 ( .A1(n317), .A2(n316), .ZN(n581) );
  AND2_X1 U438 ( .A1(a_in[0]), .A2(b_in[0]), .ZN(n579) );
  NAND2_X1 U439 ( .A1(n579), .A2(f[0]), .ZN(n584) );
  NAND2_X1 U440 ( .A1(n317), .A2(n316), .ZN(n582) );
  OAI21_X1 U441 ( .B1(n581), .B2(n584), .A(n582), .ZN(n318) );
  INV_X1 U442 ( .A(n318), .ZN(n573) );
  NAND2_X1 U443 ( .A1(n320), .A2(n319), .ZN(n571) );
  NAND2_X1 U444 ( .A1(n322), .A2(n321), .ZN(n575) );
  INV_X1 U445 ( .A(n575), .ZN(n323) );
  AOI21_X2 U446 ( .B1(n576), .B2(n577), .A(n323), .ZN(n568) );
  NAND2_X1 U447 ( .A1(n325), .A2(n324), .ZN(n566) );
  OAI21_X1 U448 ( .B1(n565), .B2(n568), .A(n566), .ZN(n556) );
  FA_X1 U449 ( .A(n327), .B(f[4]), .CI(n326), .CO(n359), .S(n336) );
  XNOR2_X1 U450 ( .A(n745), .B(a_in[0]), .ZN(n328) );
  XNOR2_X1 U451 ( .A(n745), .B(a_in[1]), .ZN(n344) );
  OAI22_X1 U452 ( .A1(n437), .A2(n328), .B1(n436), .B2(n344), .ZN(n349) );
  INV_X1 U453 ( .A(n329), .ZN(n331) );
  OR2_X1 U454 ( .A1(a_in[0]), .A2(n331), .ZN(n330) );
  OAI22_X1 U455 ( .A1(n437), .A2(n331), .B1(n330), .B2(n436), .ZN(n352) );
  XNOR2_X1 U456 ( .A(n748), .B(a_in[5]), .ZN(n355) );
  OAI22_X1 U457 ( .A1(n371), .A2(n332), .B1(n355), .B2(n765), .ZN(n351) );
  XNOR2_X1 U458 ( .A(n629), .B(a_in[3]), .ZN(n347) );
  OAI22_X1 U459 ( .A1(n348), .A2(n334), .B1(n143), .B2(n347), .ZN(n350) );
  OR2_X1 U460 ( .A1(n342), .A2(n341), .ZN(n562) );
  NAND2_X1 U461 ( .A1(n342), .A2(n341), .ZN(n561) );
  INV_X1 U462 ( .A(n561), .ZN(n555) );
  AOI21_X1 U463 ( .B1(n556), .B2(n562), .A(n555), .ZN(n388) );
  OAI22_X1 U464 ( .A1(n437), .A2(n344), .B1(n153), .B2(n343), .ZN(n362) );
  OAI22_X1 U465 ( .A1(n348), .A2(n347), .B1(n346), .B2(n345), .ZN(n361) );
  HA_X1 U466 ( .A(n349), .B(f[5]), .CO(n360), .S(n358) );
  FA_X1 U467 ( .A(n352), .B(n351), .CI(n350), .CO(n376), .S(n357) );
  INV_X1 U468 ( .A(n353), .ZN(n354) );
  AND2_X1 U469 ( .A1(a_in[0]), .A2(n354), .ZN(n368) );
  XNOR2_X1 U470 ( .A(n628), .B(a_in[6]), .ZN(n370) );
  OAI22_X1 U471 ( .A1(n371), .A2(n355), .B1(n370), .B2(n765), .ZN(n367) );
  FA_X1 U472 ( .A(n362), .B(n361), .CI(n360), .CO(n415), .S(n374) );
  FA_X1 U473 ( .A(n364), .B(n365), .CI(n363), .CO(n404), .S(n410) );
  XNOR2_X1 U474 ( .A(n415), .B(n410), .ZN(n381) );
  XNOR2_X1 U475 ( .A(n366), .B(n763), .ZN(n396) );
  FA_X1 U476 ( .A(n368), .B(f[6]), .CI(n367), .CO(n398), .S(n375) );
  OAI22_X1 U477 ( .A1(n371), .A2(n370), .B1(n369), .B2(n765), .ZN(n397) );
  XNOR2_X1 U478 ( .A(n398), .B(n397), .ZN(n372) );
  XOR2_X1 U479 ( .A(n381), .B(n414), .Z(n380) );
  INV_X1 U480 ( .A(n382), .ZN(n379) );
  NAND2_X1 U481 ( .A1(n380), .A2(n379), .ZN(n590) );
  NAND2_X1 U482 ( .A1(n558), .A2(n590), .ZN(n387) );
  XNOR2_X1 U483 ( .A(n381), .B(n414), .ZN(n383) );
  NAND2_X1 U484 ( .A1(n383), .A2(n382), .ZN(n589) );
  NAND2_X1 U485 ( .A1(n385), .A2(n384), .ZN(n559) );
  INV_X1 U486 ( .A(n559), .ZN(n587) );
  NAND2_X1 U487 ( .A1(n590), .A2(n587), .ZN(n386) );
  OAI211_X1 U488 ( .C1(n388), .C2(n387), .A(n589), .B(n386), .ZN(n546) );
  XNOR2_X1 U489 ( .A(n390), .B(n389), .ZN(n392) );
  XNOR2_X1 U490 ( .A(n392), .B(n391), .ZN(n421) );
  INV_X1 U491 ( .A(n398), .ZN(n394) );
  NAND2_X1 U492 ( .A1(n398), .A2(n397), .ZN(n399) );
  FA_X1 U493 ( .A(n403), .B(n402), .CI(n401), .CO(n233), .S(n408) );
  FA_X1 U494 ( .A(n406), .B(n405), .CI(n404), .CO(n390), .S(n407) );
  NOR2_X2 U495 ( .A1(n421), .A2(n420), .ZN(n550) );
  FA_X1 U496 ( .A(n409), .B(n408), .CI(n407), .CO(n420), .S(n419) );
  NOR2_X1 U497 ( .A1(n419), .A2(n418), .ZN(n547) );
  NOR2_X1 U498 ( .A1(n550), .A2(n547), .ZN(n423) );
  NAND2_X1 U499 ( .A1(n419), .A2(n418), .ZN(n549) );
  NAND2_X1 U500 ( .A1(n421), .A2(n420), .ZN(n551) );
  OAI21_X1 U501 ( .B1(n549), .B2(n550), .A(n551), .ZN(n422) );
  AOI21_X1 U502 ( .B1(n546), .B2(n423), .A(n422), .ZN(n504) );
  NOR2_X1 U503 ( .A1(n427), .A2(n426), .ZN(n596) );
  NAND2_X1 U504 ( .A1(n425), .A2(n424), .ZN(n606) );
  NAND2_X1 U505 ( .A1(n136), .A2(n426), .ZN(n598) );
  OAI21_X1 U506 ( .B1(n596), .B2(n606), .A(n598), .ZN(n533) );
  NAND2_X1 U507 ( .A1(n429), .A2(n428), .ZN(n537) );
  NAND2_X1 U508 ( .A1(n511), .A2(n510), .ZN(n512) );
  OAI21_X1 U509 ( .B1(n537), .B2(n152), .A(n512), .ZN(n431) );
  AOI21_X1 U510 ( .B1(n533), .B2(n432), .A(n431), .ZN(n433) );
  OAI21_X1 U511 ( .B1(n434), .B2(n137), .A(n433), .ZN(n518) );
  AOI21_X1 U512 ( .B1(n437), .B2(n153), .A(n435), .ZN(n438) );
  INV_X1 U513 ( .A(n438), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n486), .B(a_in[6]), .ZN(n449) );
  OAI22_X1 U515 ( .A1(n150), .A2(n439), .B1(n526), .B2(n449), .ZN(n452) );
  FA_X1 U516 ( .A(n441), .B(n764), .CI(n440), .CO(n451), .S(n460) );
  XNOR2_X1 U517 ( .A(n746), .B(n722), .ZN(n448) );
  OAI22_X1 U518 ( .A1(n155), .A2(n442), .B1(n471), .B2(n448), .ZN(n450) );
  OAI21_X1 U519 ( .B1(n445), .B2(n444), .A(n443), .ZN(n446) );
  NAND2_X1 U520 ( .A1(n447), .A2(n446), .ZN(n464) );
  XNOR2_X1 U521 ( .A(n746), .B(N46), .ZN(n469) );
  OAI22_X1 U522 ( .A1(n155), .A2(n448), .B1(n471), .B2(n469), .ZN(n468) );
  XNOR2_X1 U523 ( .A(a_in[7]), .B(n486), .ZN(n473) );
  OAI22_X1 U524 ( .A1(n150), .A2(n449), .B1(n526), .B2(n473), .ZN(n467) );
  FA_X1 U525 ( .A(f[13]), .B(f[14]), .CI(n450), .CO(n475), .S(n465) );
  FA_X1 U526 ( .A(n453), .B(n452), .CI(n451), .CO(n474), .S(n466) );
  NAND2_X1 U527 ( .A1(n455), .A2(n454), .ZN(n461) );
  INV_X1 U528 ( .A(n461), .ZN(n457) );
  NAND2_X1 U529 ( .A1(n457), .A2(n456), .ZN(n458) );
  FA_X1 U530 ( .A(n466), .B(n465), .CI(n464), .CO(n479), .S(n478) );
  OR2_X1 U531 ( .A1(n477), .A2(n478), .ZN(n539) );
  NAND2_X1 U532 ( .A1(n544), .A2(n539), .ZN(n499) );
  FA_X1 U533 ( .A(n468), .B(n772), .CI(n467), .CO(n491), .S(n476) );
  AOI21_X1 U534 ( .B1(n471), .B2(n154), .A(n469), .ZN(n472) );
  INV_X1 U535 ( .A(n472), .ZN(n490) );
  XNOR2_X1 U536 ( .A(n486), .B(n722), .ZN(n487) );
  OAI22_X1 U537 ( .A1(n150), .A2(n473), .B1(n526), .B2(n487), .ZN(n488) );
  FA_X1 U538 ( .A(n476), .B(n475), .CI(n474), .CO(n482), .S(n480) );
  NOR2_X1 U539 ( .A1(n483), .A2(n482), .ZN(n500) );
  NOR2_X1 U540 ( .A1(n499), .A2(n500), .ZN(n517) );
  INV_X1 U541 ( .A(n500), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n481), .A2(n544), .ZN(n485) );
  NAND2_X1 U543 ( .A1(n478), .A2(n477), .ZN(n540) );
  NAND2_X1 U544 ( .A1(n480), .A2(n479), .ZN(n543) );
  INV_X1 U545 ( .A(n543), .ZN(n496) );
  NAND2_X1 U546 ( .A1(n481), .A2(n496), .ZN(n484) );
  NAND2_X1 U547 ( .A1(n483), .A2(n482), .ZN(n501) );
  OAI211_X1 U548 ( .C1(n485), .C2(n540), .A(n484), .B(n501), .ZN(n522) );
  AOI21_X1 U549 ( .B1(n138), .B2(n517), .A(n522), .ZN(n494) );
  XNOR2_X1 U550 ( .A(n486), .B(N46), .ZN(n525) );
  OAI22_X1 U551 ( .A1(n150), .A2(n487), .B1(n526), .B2(n525), .ZN(n524) );
  FA_X1 U552 ( .A(f[15]), .B(f[16]), .CI(n488), .CO(n523), .S(n489) );
  FA_X1 U553 ( .A(n491), .B(n490), .CI(n489), .CO(n492), .S(n483) );
  OR2_X1 U554 ( .A1(n493), .A2(n492), .ZN(n521) );
  NAND2_X1 U555 ( .A1(n493), .A2(n492), .ZN(n519) );
  XNOR2_X1 U556 ( .A(n494), .B(n161), .ZN(n726) );
  INV_X1 U557 ( .A(n795), .ZN(n495) );
  INV_X1 U558 ( .A(n518), .ZN(n542) );
  OAI21_X1 U559 ( .B1(n542), .B2(n499), .A(n498), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n481), .A2(n501), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(n728) );
  INV_X1 U562 ( .A(n137), .ZN(n609) );
  INV_X1 U563 ( .A(n536), .ZN(n507) );
  NAND2_X1 U564 ( .A1(n158), .A2(n507), .ZN(n509) );
  AOI21_X1 U565 ( .B1(n534), .B2(n507), .A(n506), .ZN(n508) );
  OR2_X1 U566 ( .A1(n511), .A2(n510), .ZN(n513) );
  NAND2_X1 U567 ( .A1(n513), .A2(n512), .ZN(n514) );
  INV_X1 U568 ( .A(n519), .ZN(n520) );
  AOI21_X1 U569 ( .B1(n522), .B2(n521), .A(n520), .ZN(n614) );
  FA_X1 U570 ( .A(n524), .B(n773), .CI(n523), .CO(n529), .S(n493) );
  AOI21_X1 U571 ( .B1(n526), .B2(n150), .A(n525), .ZN(n527) );
  INV_X1 U572 ( .A(n527), .ZN(n619) );
  OR2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n615) );
  NAND2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n613) );
  NAND2_X1 U575 ( .A1(n615), .A2(n613), .ZN(n530) );
  XNOR2_X1 U576 ( .A(n531), .B(n530), .ZN(n702) );
  AND2_X1 U577 ( .A1(n540), .A2(n539), .ZN(n532) );
  XNOR2_X1 U578 ( .A(n542), .B(n532), .ZN(n680) );
  AOI21_X1 U579 ( .B1(n609), .B2(n158), .A(n534), .ZN(n538) );
  NOR2_X1 U580 ( .A1(n680), .A2(n708), .ZN(n732) );
  INV_X1 U581 ( .A(n539), .ZN(n541) );
  OAI21_X1 U582 ( .B1(n542), .B2(n541), .A(n540), .ZN(n545) );
  XNOR2_X1 U583 ( .A(n545), .B(n162), .ZN(n731) );
  INV_X1 U584 ( .A(n157), .ZN(n604) );
  INV_X1 U585 ( .A(n548), .ZN(n603) );
  OAI21_X1 U586 ( .B1(n604), .B2(n548), .A(n602), .ZN(n554) );
  INV_X1 U587 ( .A(n550), .ZN(n552) );
  NAND2_X1 U588 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U589 ( .A(n554), .B(n553), .ZN(n705) );
  AOI21_X1 U590 ( .B1(n556), .B2(n562), .A(n555), .ZN(n557) );
  INV_X1 U591 ( .A(n557), .ZN(n588) );
  NAND2_X1 U592 ( .A1(n558), .A2(n559), .ZN(n560) );
  XNOR2_X1 U593 ( .A(n588), .B(n560), .ZN(n693) );
  OAI21_X1 U594 ( .B1(n565), .B2(n568), .A(n566), .ZN(n564) );
  NAND2_X1 U595 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U596 ( .A(n564), .B(n563), .ZN(n696) );
  INV_X1 U597 ( .A(n565), .ZN(n567) );
  NAND2_X1 U598 ( .A1(n567), .A2(n566), .ZN(n569) );
  XOR2_X1 U599 ( .A(n569), .B(n568), .Z(n674) );
  INV_X1 U600 ( .A(n570), .ZN(n572) );
  NAND2_X1 U601 ( .A1(n572), .A2(n571), .ZN(n574) );
  XOR2_X1 U602 ( .A(n574), .B(n573), .Z(n638) );
  NAND2_X1 U603 ( .A1(n576), .A2(n575), .ZN(n578) );
  XNOR2_X1 U604 ( .A(n578), .B(n577), .ZN(n664) );
  OR2_X1 U605 ( .A1(n579), .A2(f[0]), .ZN(n580) );
  AND2_X1 U606 ( .A1(n580), .A2(n584), .ZN(n661) );
  INV_X1 U607 ( .A(n581), .ZN(n583) );
  NAND2_X1 U608 ( .A1(n583), .A2(n582), .ZN(n585) );
  XOR2_X1 U609 ( .A(n585), .B(n584), .Z(n671) );
  OR4_X1 U610 ( .A1(n638), .A2(n664), .A3(n661), .A4(n671), .ZN(n586) );
  OR4_X1 U611 ( .A1(n693), .A2(n696), .A3(n674), .A4(n586), .ZN(n593) );
  AOI21_X1 U612 ( .B1(n588), .B2(n558), .A(n587), .ZN(n592) );
  NAND2_X1 U613 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U614 ( .A(n592), .B(n591), .Z(n699) );
  OR3_X1 U615 ( .A1(n705), .A2(n593), .A3(n699), .ZN(n610) );
  INV_X1 U616 ( .A(n594), .ZN(n607) );
  INV_X1 U617 ( .A(n606), .ZN(n595) );
  AOI21_X1 U618 ( .B1(n609), .B2(n607), .A(n595), .ZN(n601) );
  INV_X1 U619 ( .A(n597), .ZN(n599) );
  NAND2_X1 U620 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U621 ( .A(n601), .B(n600), .Z(n686) );
  NAND2_X1 U622 ( .A1(n603), .A2(n602), .ZN(n605) );
  XOR2_X1 U623 ( .A(n605), .B(n604), .Z(n683) );
  NAND2_X1 U624 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U625 ( .A(n609), .B(n608), .ZN(n677) );
  NOR4_X2 U626 ( .A1(n610), .A2(n686), .A3(n683), .A4(n677), .ZN(n730) );
  NAND3_X1 U627 ( .A1(n612), .A2(n611), .A3(n730), .ZN(n660) );
  AND2_X1 U628 ( .A1(n614), .A2(n613), .ZN(n618) );
  INV_X1 U629 ( .A(n615), .ZN(n616) );
  FA_X1 U630 ( .A(f[17]), .B(f[18]), .CI(n619), .CO(n620), .S(n528) );
  OR2_X1 U631 ( .A1(n620), .A2(n769), .ZN(n622) );
  NAND2_X1 U632 ( .A1(n620), .A2(n769), .ZN(n621) );
  NOR3_X1 U633 ( .A1(a_in[0]), .A2(a_in[7]), .A3(n722), .ZN(n627) );
  NOR2_X1 U634 ( .A1(a_in[5]), .A2(a_in[6]), .ZN(n626) );
  NOR2_X1 U635 ( .A1(a_in[3]), .A2(a_in[4]), .ZN(n625) );
  NOR2_X1 U636 ( .A1(a_in[2]), .A2(a_in[1]), .ZN(n624) );
  NAND4_X1 U637 ( .A1(n627), .A2(n626), .A3(n625), .A4(n624), .ZN(n639) );
  AND2_X1 U638 ( .A1(n639), .A2(n486), .ZN(n636) );
  NOR3_X1 U639 ( .A1(n628), .A2(b_in[6]), .A3(b_in[4]), .ZN(n633) );
  NOR2_X1 U640 ( .A1(b_in[8]), .A2(b_in[2]), .ZN(n632) );
  NOR2_X1 U641 ( .A1(n746), .A2(b_in[0]), .ZN(n631) );
  NOR2_X1 U642 ( .A1(n745), .A2(n743), .ZN(n630) );
  NAND4_X1 U643 ( .A1(n633), .A2(n632), .A3(n631), .A4(n630), .ZN(n634) );
  NAND2_X1 U644 ( .A1(n634), .A2(n766), .ZN(n641) );
  NAND2_X1 U645 ( .A1(n641), .A2(N46), .ZN(n635) );
  OAI211_X1 U646 ( .C1(n636), .C2(N46), .A(N55), .B(n635), .ZN(n637) );
  OR2_X1 U647 ( .A1(n735), .A2(n637), .ZN(n734) );
  NAND2_X1 U648 ( .A1(n734), .A2(n795), .ZN(n659) );
  NAND2_X1 U649 ( .A1(n660), .A2(n659), .ZN(n712) );
  NAND2_X1 U650 ( .A1(n712), .A2(n638), .ZN(n658) );
  INV_X1 U651 ( .A(n639), .ZN(n640) );
  OR2_X1 U652 ( .A1(n641), .A2(n640), .ZN(n655) );
  OR2_X1 U653 ( .A1(f[18]), .A2(f[1]), .ZN(n642) );
  NOR3_X1 U654 ( .A1(n642), .A2(f[5]), .A3(f[3]), .ZN(n646) );
  NOR3_X1 U655 ( .A1(f[0]), .A2(f[9]), .A3(f[7]), .ZN(n645) );
  NOR2_X1 U656 ( .A1(f[15]), .A2(f[13]), .ZN(n644) );
  NOR2_X1 U657 ( .A1(f[10]), .A2(f[11]), .ZN(n643) );
  NAND4_X1 U658 ( .A1(n646), .A2(n645), .A3(n644), .A4(n643), .ZN(n653) );
  NOR2_X1 U659 ( .A1(f[16]), .A2(f[14]), .ZN(n650) );
  NOR2_X1 U660 ( .A1(f[12]), .A2(f[8]), .ZN(n649) );
  NOR2_X1 U661 ( .A1(f[6]), .A2(f[4]), .ZN(n648) );
  NOR2_X1 U662 ( .A1(f[17]), .A2(f[2]), .ZN(n647) );
  NAND4_X1 U663 ( .A1(n650), .A2(n649), .A3(n648), .A4(n647), .ZN(n652) );
  AOI21_X1 U664 ( .B1(n766), .B2(N46), .A(N55), .ZN(n651) );
  OAI21_X1 U665 ( .B1(n653), .B2(n652), .A(n651), .ZN(n654) );
  AOI21_X1 U666 ( .B1(n752), .B2(n655), .A(n654), .ZN(n656) );
  AND2_X2 U667 ( .A1(n735), .A2(n656), .ZN(n738) );
  NAND2_X2 U668 ( .A1(n738), .A2(n795), .ZN(n713) );
  INV_X1 U669 ( .A(reset), .ZN(n716) );
  AND2_X1 U670 ( .A1(n713), .A2(n166), .ZN(n657) );
  NAND2_X1 U671 ( .A1(n658), .A2(n657), .ZN(n95) );
  NAND2_X1 U672 ( .A1(n712), .A2(n661), .ZN(n663) );
  AND2_X1 U673 ( .A1(n713), .A2(n167), .ZN(n662) );
  NAND2_X1 U674 ( .A1(n663), .A2(n662), .ZN(n97) );
  NAND2_X1 U675 ( .A1(n147), .A2(n664), .ZN(n666) );
  AND2_X1 U676 ( .A1(n713), .A2(n168), .ZN(n665) );
  NAND2_X1 U677 ( .A1(n666), .A2(n665), .ZN(n94) );
  INV_X1 U678 ( .A(n667), .ZN(n668) );
  NAND2_X1 U679 ( .A1(n148), .A2(n668), .ZN(n670) );
  AND2_X1 U680 ( .A1(n713), .A2(n169), .ZN(n669) );
  NAND2_X1 U681 ( .A1(n670), .A2(n669), .ZN(n82) );
  NAND2_X1 U682 ( .A1(n709), .A2(n671), .ZN(n673) );
  AND2_X1 U683 ( .A1(n713), .A2(n170), .ZN(n672) );
  NAND2_X1 U684 ( .A1(n673), .A2(n672), .ZN(n96) );
  NAND2_X1 U685 ( .A1(n147), .A2(n674), .ZN(n676) );
  AND2_X1 U686 ( .A1(n713), .A2(n171), .ZN(n675) );
  NAND2_X1 U687 ( .A1(n676), .A2(n675), .ZN(n93) );
  NAND2_X1 U688 ( .A1(n709), .A2(n677), .ZN(n679) );
  AND2_X1 U689 ( .A1(n713), .A2(n172), .ZN(n678) );
  NAND2_X1 U690 ( .A1(n679), .A2(n678), .ZN(n87) );
  NAND2_X1 U691 ( .A1(n148), .A2(n680), .ZN(n682) );
  AND2_X1 U692 ( .A1(n713), .A2(n173), .ZN(n681) );
  NAND2_X1 U693 ( .A1(n682), .A2(n681), .ZN(n83) );
  NAND2_X1 U694 ( .A1(n147), .A2(n683), .ZN(n685) );
  AND2_X1 U695 ( .A1(n713), .A2(n174), .ZN(n684) );
  NAND2_X1 U696 ( .A1(n685), .A2(n684), .ZN(n89) );
  NAND2_X1 U697 ( .A1(n712), .A2(n686), .ZN(n688) );
  AND2_X1 U698 ( .A1(n713), .A2(n175), .ZN(n687) );
  NAND2_X1 U699 ( .A1(n688), .A2(n687), .ZN(n86) );
  NAND2_X1 U700 ( .A1(n709), .A2(n142), .ZN(n690) );
  AND2_X1 U701 ( .A1(n713), .A2(n176), .ZN(n689) );
  NAND2_X1 U702 ( .A1(n690), .A2(n689), .ZN(n80) );
  NAND2_X1 U703 ( .A1(n148), .A2(n156), .ZN(n692) );
  AND2_X1 U704 ( .A1(n713), .A2(n177), .ZN(n691) );
  NAND2_X1 U705 ( .A1(n692), .A2(n691), .ZN(n81) );
  NAND2_X1 U706 ( .A1(n712), .A2(n693), .ZN(n695) );
  NAND2_X1 U707 ( .A1(n695), .A2(n694), .ZN(n91) );
  NAND2_X1 U708 ( .A1(n147), .A2(n696), .ZN(n698) );
  NAND2_X1 U709 ( .A1(n698), .A2(n697), .ZN(n92) );
  NAND2_X1 U710 ( .A1(n148), .A2(n699), .ZN(n701) );
  NAND2_X1 U711 ( .A1(n701), .A2(n700), .ZN(n90) );
  NAND2_X1 U712 ( .A1(n712), .A2(n702), .ZN(n704) );
  NAND2_X1 U713 ( .A1(n704), .A2(n703), .ZN(n79) );
  NAND2_X1 U714 ( .A1(n147), .A2(n705), .ZN(n707) );
  AND2_X1 U715 ( .A1(n713), .A2(n178), .ZN(n706) );
  NAND2_X1 U716 ( .A1(n707), .A2(n706), .ZN(n88) );
  NAND2_X1 U717 ( .A1(n709), .A2(n708), .ZN(n711) );
  AND2_X1 U718 ( .A1(n713), .A2(n179), .ZN(n710) );
  NAND2_X1 U719 ( .A1(n711), .A2(n710), .ZN(n85) );
  NAND2_X1 U720 ( .A1(n148), .A2(n727), .ZN(n715) );
  AND2_X1 U721 ( .A1(n713), .A2(n180), .ZN(n714) );
  NAND2_X1 U722 ( .A1(n715), .A2(n714), .ZN(n84) );
  NOR2_X2 U723 ( .A1(valid_in), .A2(reset), .ZN(n749) );
  AOI22_X1 U724 ( .A1(n796), .A2(a[0]), .B1(n749), .B2(a_in[0]), .ZN(n790) );
  AOI22_X1 U725 ( .A1(n796), .A2(b[6]), .B1(n749), .B2(b_in[6]), .ZN(n792) );
  AOI22_X1 U726 ( .A1(n796), .A2(b[8]), .B1(n749), .B2(b_in[8]), .ZN(n717) );
  INV_X1 U727 ( .A(n717), .ZN(n106) );
  AOI22_X1 U728 ( .A1(n796), .A2(b[0]), .B1(n749), .B2(b_in[0]), .ZN(n794) );
  AOI22_X1 U729 ( .A1(n796), .A2(b[2]), .B1(n749), .B2(b_in[2]), .ZN(n793) );
  AOI22_X1 U730 ( .A1(n796), .A2(a[2]), .B1(n749), .B2(a_in[2]), .ZN(n789) );
  AOI22_X1 U731 ( .A1(n796), .A2(a[3]), .B1(n749), .B2(a_in[3]), .ZN(n788) );
  AOI22_X1 U732 ( .A1(n796), .A2(a[4]), .B1(n749), .B2(a_in[4]), .ZN(n718) );
  INV_X1 U733 ( .A(n718), .ZN(n112) );
  AOI22_X1 U734 ( .A1(n796), .A2(a[5]), .B1(n749), .B2(a_in[5]), .ZN(n719) );
  INV_X1 U735 ( .A(n719), .ZN(n113) );
  AOI22_X1 U736 ( .A1(n796), .A2(a[1]), .B1(n749), .B2(a_in[1]), .ZN(n720) );
  INV_X1 U737 ( .A(n720), .ZN(n109) );
  AOI22_X1 U738 ( .A1(n796), .A2(a[7]), .B1(n749), .B2(a_in[7]), .ZN(n721) );
  INV_X1 U739 ( .A(n721), .ZN(n115) );
  AOI22_X1 U740 ( .A1(n796), .A2(a[8]), .B1(n749), .B2(n722), .ZN(n723) );
  INV_X1 U741 ( .A(n723), .ZN(n116) );
  AOI22_X1 U742 ( .A1(n796), .A2(a[9]), .B1(n749), .B2(N46), .ZN(n724) );
  INV_X1 U743 ( .A(n724), .ZN(n117) );
  AOI22_X1 U744 ( .A1(n796), .A2(b[4]), .B1(n749), .B2(b_in[4]), .ZN(n725) );
  INV_X1 U745 ( .A(n725), .ZN(n102) );
  AOI22_X1 U746 ( .A1(n796), .A2(a[6]), .B1(n749), .B2(a_in[6]), .ZN(n787) );
  NOR3_X1 U747 ( .A1(n134), .A2(n727), .A3(n142), .ZN(n729) );
  AND2_X1 U748 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U749 ( .A1(n733), .A2(n611), .ZN(n737) );
  INV_X1 U750 ( .A(n734), .ZN(n736) );
  AOI21_X1 U751 ( .B1(n737), .B2(n736), .A(n735), .ZN(n742) );
  INV_X1 U752 ( .A(n738), .ZN(n739) );
  NAND2_X1 U753 ( .A1(n739), .A2(n795), .ZN(n741) );
  OAI22_X1 U754 ( .A1(n742), .A2(n741), .B1(n740), .B2(n769), .ZN(n78) );
  AOI22_X1 U755 ( .A1(n796), .A2(b[3]), .B1(n749), .B2(n743), .ZN(n744) );
  INV_X1 U756 ( .A(n744), .ZN(n101) );
  AOI22_X1 U757 ( .A1(n796), .A2(b[5]), .B1(n749), .B2(n745), .ZN(n785) );
  AOI22_X1 U758 ( .A1(n796), .A2(b[7]), .B1(n749), .B2(n746), .ZN(n747) );
  INV_X1 U759 ( .A(n747), .ZN(n105) );
  AOI22_X1 U760 ( .A1(n796), .A2(b[1]), .B1(n749), .B2(n748), .ZN(n786) );
  AOI22_X1 U761 ( .A1(n796), .A2(b[9]), .B1(n749), .B2(n486), .ZN(n791) );
endmodule

