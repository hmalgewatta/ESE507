
module part1_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   enable_f, n47, n48, n49, n50, n51, n52, n53, n54, n56, n57, n60, n61,
         n62, n63, n64, n65, n66, n67, n70, n72, n73, n77, n78, n79, n80, n81,
         n83, n84, n85, n86, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665;
  wire   [9:0] a_in;
  wire   [9:0] b_in;

  DFF_X1 \f_reg[14]  ( .D(n53), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[13]  ( .D(n54), .CK(clk), .Q(f[13]), .QN(n146) );
  DFF_X1 \f_reg[12]  ( .D(n638), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[11]  ( .D(n56), .CK(clk), .Q(f[11]), .QN(n145) );
  DFF_X1 \f_reg[10]  ( .D(n57), .CK(clk), .Q(f[10]) );
  DFF_X1 \a_in_reg[9]  ( .D(n77), .CK(clk), .Q(a_in[9]) );
  DFF_X1 \a_in_reg[8]  ( .D(n78), .CK(clk), .Q(a_in[8]) );
  DFF_X1 \a_in_reg[7]  ( .D(n79), .CK(clk), .Q(a_in[7]) );
  DFF_X1 \a_in_reg[6]  ( .D(n80), .CK(clk), .Q(a_in[6]) );
  DFF_X1 \a_in_reg[5]  ( .D(n81), .CK(clk), .Q(a_in[5]) );
  DFF_X1 \a_in_reg[3]  ( .D(n83), .CK(clk), .Q(a_in[3]) );
  DFF_X1 \a_in_reg[2]  ( .D(n84), .CK(clk), .Q(a_in[2]) );
  DFF_X1 \a_in_reg[1]  ( .D(n85), .CK(clk), .Q(a_in[1]) );
  DFF_X1 \b_in_reg[4]  ( .D(n73), .CK(clk), .Q(b_in[4]), .QN(n642) );
  DFF_X1 \b_in_reg[7]  ( .D(n70), .CK(clk), .Q(b_in[7]), .QN(n663) );
  DFF_X1 \f_reg[19]  ( .D(n48), .CK(clk), .Q(f[19]), .QN(n648) );
  DFF_X1 \b_in_reg[9]  ( .D(n654), .CK(clk), .Q(n641), .QN(b_in[9]) );
  DFF_X1 \b_in_reg[8]  ( .D(n657), .CK(clk), .Q(n640), .QN(b_in[8]) );
  DFF_X1 \b_in_reg[3]  ( .D(n655), .CK(clk), .Q(n643), .QN(b_in[3]) );
  DFF_X1 \b_in_reg[2]  ( .D(n659), .CK(clk), .Q(n647), .QN(b_in[2]) );
  DFF_X1 \b_in_reg[1]  ( .D(n653), .CK(clk), .Q(n644), .QN(b_in[1]) );
  DFF_X2 \f_reg[16]  ( .D(n51), .CK(clk), .Q(f[16]) );
  DFF_X2 \f_reg[18]  ( .D(n49), .CK(clk), .Q(f[18]) );
  DFF_X2 \f_reg[15]  ( .D(n52), .CK(clk), .Q(f[15]), .QN(n650) );
  DFF_X2 \f_reg[17]  ( .D(n50), .CK(clk), .Q(f[17]), .QN(n649) );
  DFF_X1 valid_out_reg ( .D(n665), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[0]  ( .D(n67), .CK(clk), .Q(f[0]) );
  DFF_X1 \f_reg[1]  ( .D(n66), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[2]  ( .D(n65), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(n64), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(n63), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(n62), .CK(clk), .Q(f[5]), .QN(n102) );
  DFF_X1 \f_reg[6]  ( .D(n61), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(n60), .CK(clk), .Q(f[7]), .QN(n645) );
  DFF_X1 \f_reg[8]  ( .D(n662), .CK(clk), .QN(f[8]) );
  DFF_X1 \f_reg[9]  ( .D(n661), .CK(clk), .Q(n646), .QN(f[9]) );
  DFF_X1 \a_in_reg[4]  ( .D(n656), .CK(clk), .QN(a_in[4]) );
  SDFF_X1 enable_f_reg ( .D(n47), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(enable_f), 
        .QN(n652) );
  DFF_X1 \b_in_reg[0]  ( .D(n660), .CK(clk), .Q(n651), .QN(b_in[0]) );
  DFF_X1 \b_in_reg[6]  ( .D(n658), .CK(clk), .Q(n639), .QN(b_in[6]) );
  DFF_X2 \a_in_reg[0]  ( .D(n86), .CK(clk), .Q(a_in[0]), .QN(n144) );
  DFF_X1 \b_in_reg[5]  ( .D(n72), .CK(clk), .Q(b_in[5]), .QN(n664) );
  XNOR2_X1 U91 ( .A(n95), .B(n96), .ZN(n311) );
  NAND2_X1 U92 ( .A1(n460), .A2(n461), .ZN(n98) );
  XNOR2_X1 U93 ( .A(n309), .B(n308), .ZN(n96) );
  OR2_X1 U94 ( .A1(n435), .A2(n449), .ZN(n92) );
  XNOR2_X1 U95 ( .A(n91), .B(n90), .ZN(n228) );
  OR2_X1 U96 ( .A1(n242), .A2(n358), .ZN(n245) );
  XNOR2_X1 U97 ( .A(n219), .B(f[6]), .ZN(n91) );
  INV_X1 U98 ( .A(n386), .ZN(n426) );
  OR2_X1 U99 ( .A1(n644), .A2(b_in[0]), .ZN(n299) );
  NAND2_X2 U100 ( .A1(n190), .A2(n189), .ZN(n193) );
  INV_X2 U101 ( .A(n663), .ZN(n431) );
  NAND2_X1 U102 ( .A1(n89), .A2(n88), .ZN(n241) );
  NAND2_X2 U103 ( .A1(n90), .A2(f[6]), .ZN(n88) );
  OAI21_X2 U104 ( .B1(n90), .B2(f[6]), .A(n219), .ZN(n89) );
  OAI22_X2 U105 ( .A1(n203), .A2(n651), .B1(n202), .B2(n299), .ZN(n90) );
  NOR2_X1 U106 ( .A1(n414), .A2(n413), .ZN(n419) );
  NOR2_X1 U107 ( .A1(n407), .A2(n406), .ZN(n414) );
  OAI21_X1 U108 ( .B1(n293), .B2(n292), .A(n291), .ZN(n116) );
  NOR2_X1 U109 ( .A1(n338), .A2(n339), .ZN(n413) );
  OAI21_X2 U110 ( .B1(n450), .B2(n392), .A(n92), .ZN(n466) );
  AOI21_X1 U111 ( .B1(n603), .B2(n290), .A(n289), .ZN(n138) );
  OAI21_X1 U112 ( .B1(n610), .B2(n607), .A(n611), .ZN(n289) );
  NAND2_X1 U113 ( .A1(n235), .A2(n234), .ZN(n596) );
  XNOR2_X1 U114 ( .A(n258), .B(n217), .ZN(n235) );
  NAND2_X1 U115 ( .A1(n94), .A2(n93), .ZN(n315) );
  NAND2_X1 U116 ( .A1(n309), .A2(n308), .ZN(n93) );
  OAI21_X1 U117 ( .B1(n308), .B2(n309), .A(n95), .ZN(n94) );
  XNOR2_X1 U118 ( .A(n296), .B(n646), .ZN(n95) );
  NAND2_X1 U119 ( .A1(n97), .A2(n501), .ZN(n508) );
  AND2_X1 U120 ( .A1(n498), .A2(n665), .ZN(n97) );
  AOI21_X2 U121 ( .B1(n622), .B2(n536), .A(n487), .ZN(n527) );
  NAND2_X2 U122 ( .A1(n99), .A2(n98), .ZN(n472) );
  NAND2_X2 U123 ( .A1(n459), .A2(n100), .ZN(n99) );
  OR2_X2 U124 ( .A1(n460), .A2(n461), .ZN(n100) );
  XNOR2_X1 U125 ( .A(n101), .B(n459), .ZN(n477) );
  XNOR2_X1 U126 ( .A(n460), .B(n461), .ZN(n101) );
  NAND2_X1 U127 ( .A1(n293), .A2(n292), .ZN(n115) );
  NAND2_X1 U128 ( .A1(n369), .A2(n368), .ZN(n118) );
  XNOR2_X1 U129 ( .A(n369), .B(n368), .ZN(n128) );
  AOI21_X1 U130 ( .B1(n193), .B2(n105), .A(n664), .ZN(n222) );
  BUF_X2 U131 ( .A(n160), .Z(n362) );
  BUF_X1 U132 ( .A(b_in[9]), .Z(n136) );
  BUF_X1 U133 ( .A(b_in[1]), .Z(n248) );
  NAND2_X1 U134 ( .A1(n372), .A2(n421), .ZN(n373) );
  INV_X1 U135 ( .A(n414), .ZN(n137) );
  INV_X1 U136 ( .A(n413), .ZN(n141) );
  BUF_X1 U137 ( .A(n418), .Z(n378) );
  NAND2_X1 U138 ( .A1(n132), .A2(n131), .ZN(n339) );
  NAND2_X1 U139 ( .A1(n337), .A2(n336), .ZN(n131) );
  NAND2_X1 U140 ( .A1(n122), .A2(n121), .ZN(n483) );
  NAND2_X1 U141 ( .A1(n471), .A2(n470), .ZN(n121) );
  XNOR2_X1 U142 ( .A(n114), .B(n113), .ZN(n286) );
  NAND2_X1 U143 ( .A1(n116), .A2(n115), .ZN(n337) );
  OAI21_X1 U144 ( .B1(n471), .B2(n470), .A(n469), .ZN(n122) );
  NAND2_X1 U145 ( .A1(n125), .A2(n124), .ZN(n234) );
  XNOR2_X1 U146 ( .A(n284), .B(n283), .ZN(n114) );
  OR2_X1 U147 ( .A1(n233), .A2(n232), .ZN(n594) );
  NAND2_X1 U148 ( .A1(n108), .A2(n107), .ZN(n185) );
  NAND2_X1 U149 ( .A1(n226), .A2(n126), .ZN(n125) );
  XNOR2_X1 U150 ( .A(n228), .B(n227), .ZN(n127) );
  OR2_X1 U151 ( .A1(n227), .A2(n228), .ZN(n126) );
  NAND2_X1 U152 ( .A1(n274), .A2(n275), .ZN(n276) );
  NAND2_X1 U153 ( .A1(n228), .A2(n227), .ZN(n124) );
  NAND2_X1 U154 ( .A1(n167), .A2(n109), .ZN(n108) );
  NAND2_X1 U155 ( .A1(n317), .A2(n316), .ZN(n129) );
  OR2_X1 U156 ( .A1(n169), .A2(n168), .ZN(n109) );
  AND2_X1 U157 ( .A1(n216), .A2(f[5]), .ZN(n223) );
  NAND2_X1 U158 ( .A1(n169), .A2(n168), .ZN(n107) );
  BUF_X1 U159 ( .A(n348), .Z(n142) );
  NAND2_X1 U160 ( .A1(n211), .A2(n144), .ZN(n105) );
  INV_X1 U161 ( .A(n211), .ZN(n359) );
  INV_X1 U162 ( .A(n206), .ZN(n435) );
  BUF_X2 U163 ( .A(b_in[9]), .Z(n631) );
  AND2_X1 U164 ( .A1(valid_in), .A2(n540), .ZN(n635) );
  AOI21_X1 U165 ( .B1(n651), .B2(n299), .A(n298), .ZN(n300) );
  XNOR2_X1 U166 ( .A(a_in[9]), .B(b_in[1]), .ZN(n298) );
  NAND2_X1 U167 ( .A1(n233), .A2(n232), .ZN(n589) );
  XNOR2_X1 U168 ( .A(n127), .B(n226), .ZN(n233) );
  XNOR2_X1 U169 ( .A(n104), .B(n147), .ZN(n405) );
  NAND2_X1 U170 ( .A1(n381), .A2(n382), .ZN(n104) );
  OAI21_X1 U171 ( .B1(n106), .B2(n499), .A(n375), .ZN(n638) );
  XNOR2_X1 U172 ( .A(n374), .B(n373), .ZN(n106) );
  OR2_X2 U173 ( .A1(n235), .A2(n234), .ZN(n597) );
  OAI21_X1 U174 ( .B1(n337), .B2(n336), .A(n133), .ZN(n132) );
  XNOR2_X1 U175 ( .A(n167), .B(n110), .ZN(n183) );
  XNOR2_X1 U176 ( .A(n169), .B(n168), .ZN(n110) );
  NAND2_X1 U177 ( .A1(n112), .A2(n111), .ZN(n287) );
  NAND2_X1 U178 ( .A1(n284), .A2(n283), .ZN(n111) );
  OAI21_X1 U179 ( .B1(n283), .B2(n284), .A(n113), .ZN(n112) );
  XNOR2_X1 U180 ( .A(n254), .B(n273), .ZN(n113) );
  XNOR2_X1 U181 ( .A(n469), .B(n470), .ZN(n123) );
  XNOR2_X1 U182 ( .A(n394), .B(n464), .ZN(n469) );
  XNOR2_X1 U183 ( .A(n117), .B(n291), .ZN(n310) );
  XNOR2_X1 U184 ( .A(n293), .B(n292), .ZN(n117) );
  OAI21_X1 U185 ( .B1(n369), .B2(n368), .A(n367), .ZN(n119) );
  NAND2_X1 U186 ( .A1(n119), .A2(n118), .ZN(n370) );
  AOI21_X1 U187 ( .B1(n583), .B2(n585), .A(n201), .ZN(n588) );
  OAI21_X1 U188 ( .B1(n578), .B2(n575), .A(n576), .ZN(n585) );
  NAND2_X2 U189 ( .A1(n130), .A2(n129), .ZN(n369) );
  XNOR2_X1 U190 ( .A(n331), .B(n332), .ZN(n297) );
  XNOR2_X1 U191 ( .A(n320), .B(f[10]), .ZN(n331) );
  NAND2_X1 U192 ( .A1(n286), .A2(n285), .ZN(n607) );
  BUF_X4 U193 ( .A(b_in[3]), .Z(n633) );
  OAI21_X1 U194 ( .B1(n316), .B2(n317), .A(n315), .ZN(n130) );
  NOR2_X1 U195 ( .A1(n339), .A2(n340), .ZN(n342) );
  XNOR2_X1 U196 ( .A(n120), .B(n367), .ZN(n340) );
  XNOR2_X1 U197 ( .A(n369), .B(n368), .ZN(n120) );
  OAI21_X1 U198 ( .B1(n588), .B2(n238), .A(n237), .ZN(n139) );
  AOI21_X1 U199 ( .B1(n593), .B2(n597), .A(n236), .ZN(n237) );
  XNOR2_X1 U200 ( .A(n216), .B(n102), .ZN(n230) );
  XNOR2_X1 U201 ( .A(n123), .B(n471), .ZN(n416) );
  XNOR2_X1 U202 ( .A(n128), .B(n367), .ZN(n338) );
  XNOR2_X1 U203 ( .A(n135), .B(n133), .ZN(n407) );
  XNOR2_X1 U204 ( .A(n315), .B(n134), .ZN(n133) );
  XNOR2_X1 U205 ( .A(n317), .B(n316), .ZN(n134) );
  XNOR2_X1 U206 ( .A(n337), .B(n336), .ZN(n135) );
  AOI21_X1 U207 ( .B1(n139), .B2(n290), .A(n289), .ZN(n511) );
  NAND2_X1 U208 ( .A1(n205), .A2(n204), .ZN(n140) );
  NAND2_X1 U209 ( .A1(n205), .A2(n204), .ZN(n358) );
  OAI22_X1 U210 ( .A1(n445), .A2(n322), .B1(n143), .B2(n346), .ZN(n348) );
  BUF_X1 U211 ( .A(n321), .Z(n143) );
  AND2_X1 U212 ( .A1(f[9]), .A2(n296), .ZN(n333) );
  NAND2_X1 U213 ( .A1(n350), .A2(n349), .ZN(n384) );
  NAND2_X1 U214 ( .A1(n333), .A2(n332), .ZN(n334) );
  NAND2_X1 U215 ( .A1(n328), .A2(n327), .ZN(n329) );
  INV_X1 U216 ( .A(n259), .ZN(n255) );
  XNOR2_X1 U217 ( .A(n250), .B(n645), .ZN(n239) );
  XNOR2_X1 U218 ( .A(n647), .B(b_in[3]), .ZN(n159) );
  XNOR2_X1 U219 ( .A(n297), .B(n333), .ZN(n336) );
  NAND2_X1 U220 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U221 ( .A(b_in[1]), .B(b_in[2]), .ZN(n160) );
  NAND2_X1 U222 ( .A1(n310), .A2(n153), .ZN(n314) );
  NAND2_X1 U223 ( .A1(n330), .A2(n329), .ZN(n355) );
  NAND2_X1 U224 ( .A1(n262), .A2(n261), .ZN(n285) );
  NAND2_X1 U225 ( .A1(n258), .A2(n257), .ZN(n262) );
  NAND2_X1 U226 ( .A1(n256), .A2(n255), .ZN(n257) );
  NAND2_X1 U227 ( .A1(n468), .A2(n467), .ZN(n475) );
  NAND2_X1 U228 ( .A1(n464), .A2(n463), .ZN(n468) );
  OAI21_X1 U229 ( .B1(n412), .B2(n499), .A(n411), .ZN(n56) );
  NAND2_X1 U230 ( .A1(n627), .A2(f[11]), .ZN(n411) );
  AND2_X1 U231 ( .A1(enable_f), .A2(n540), .ZN(n665) );
  AND2_X1 U232 ( .A1(n403), .A2(n420), .ZN(n147) );
  NAND2_X1 U233 ( .A1(n521), .A2(n525), .ZN(n148) );
  NAND2_X1 U234 ( .A1(n516), .A2(n515), .ZN(n149) );
  NAND2_X1 U235 ( .A1(n531), .A2(n530), .ZN(n150) );
  NAND2_X1 U236 ( .A1(n536), .A2(n535), .ZN(n151) );
  AND2_X1 U237 ( .A1(n502), .A2(n503), .ZN(n152) );
  OR2_X1 U238 ( .A1(n312), .A2(n311), .ZN(n153) );
  NAND2_X1 U239 ( .A1(n627), .A2(f[18]), .ZN(n154) );
  NAND2_X1 U240 ( .A1(n627), .A2(f[16]), .ZN(n155) );
  NAND2_X1 U241 ( .A1(n627), .A2(f[17]), .ZN(n156) );
  NAND2_X1 U242 ( .A1(n627), .A2(f[15]), .ZN(n157) );
  OR2_X1 U243 ( .A1(n498), .A2(n505), .ZN(n158) );
  XNOR2_X1 U245 ( .A(n248), .B(a_in[2]), .ZN(n171) );
  XNOR2_X1 U246 ( .A(n248), .B(a_in[3]), .ZN(n161) );
  OAI22_X1 U247 ( .A1(n299), .A2(n171), .B1(n161), .B2(n651), .ZN(n166) );
  NAND2_X2 U248 ( .A1(n160), .A2(n159), .ZN(n361) );
  XNOR2_X1 U249 ( .A(n633), .B(a_in[1]), .ZN(n164) );
  XNOR2_X1 U250 ( .A(n633), .B(a_in[2]), .ZN(n195) );
  OAI22_X1 U251 ( .A1(n361), .A2(n164), .B1(n362), .B2(n195), .ZN(n197) );
  XNOR2_X1 U252 ( .A(n642), .B(n643), .ZN(n189) );
  INV_X1 U253 ( .A(n189), .ZN(n211) );
  AND2_X1 U254 ( .A1(n211), .A2(a_in[0]), .ZN(n188) );
  INV_X1 U255 ( .A(n644), .ZN(n630) );
  XNOR2_X1 U256 ( .A(n630), .B(a_in[4]), .ZN(n194) );
  OAI22_X1 U257 ( .A1(n299), .A2(n161), .B1(n194), .B2(n651), .ZN(n187) );
  INV_X1 U258 ( .A(n633), .ZN(n163) );
  OR2_X1 U259 ( .A1(a_in[0]), .A2(n163), .ZN(n162) );
  OAI22_X1 U260 ( .A1(n361), .A2(n163), .B1(n162), .B2(n362), .ZN(n169) );
  XNOR2_X1 U261 ( .A(n633), .B(a_in[0]), .ZN(n165) );
  OAI22_X1 U262 ( .A1(n361), .A2(n165), .B1(n362), .B2(n164), .ZN(n168) );
  HA_X1 U263 ( .A(n166), .B(f[3]), .CO(n198), .S(n167) );
  NOR2_X1 U264 ( .A1(n186), .A2(n185), .ZN(n575) );
  INV_X1 U265 ( .A(n362), .ZN(n170) );
  AND2_X1 U266 ( .A1(a_in[0]), .A2(n170), .ZN(n173) );
  XNOR2_X1 U267 ( .A(n630), .B(a_in[1]), .ZN(n174) );
  OAI22_X1 U268 ( .A1(n299), .A2(n174), .B1(n171), .B2(n651), .ZN(n172) );
  OR2_X1 U269 ( .A1(n183), .A2(n182), .ZN(n563) );
  FA_X1 U270 ( .A(n172), .B(f[2]), .CI(n173), .CO(n182), .S(n181) );
  OAI22_X1 U271 ( .A1(n299), .A2(a_in[0]), .B1(n174), .B2(n651), .ZN(n175) );
  NOR2_X1 U272 ( .A1(n181), .A2(n180), .ZN(n568) );
  HA_X1 U273 ( .A(n175), .B(f[1]), .CO(n180), .S(n178) );
  OR2_X1 U274 ( .A1(a_in[0]), .A2(n644), .ZN(n176) );
  NAND2_X1 U275 ( .A1(n176), .A2(n299), .ZN(n177) );
  NOR2_X1 U276 ( .A1(n178), .A2(n177), .ZN(n555) );
  AND2_X1 U277 ( .A1(a_in[0]), .A2(b_in[0]), .ZN(n541) );
  NAND2_X1 U278 ( .A1(n541), .A2(f[0]), .ZN(n558) );
  NAND2_X1 U279 ( .A1(n178), .A2(n177), .ZN(n556) );
  OAI21_X1 U280 ( .B1(n555), .B2(n558), .A(n556), .ZN(n179) );
  INV_X1 U281 ( .A(n179), .ZN(n571) );
  NAND2_X1 U282 ( .A1(n181), .A2(n180), .ZN(n569) );
  OAI21_X1 U283 ( .B1(n568), .B2(n571), .A(n569), .ZN(n564) );
  NAND2_X1 U284 ( .A1(n183), .A2(n182), .ZN(n562) );
  INV_X1 U285 ( .A(n562), .ZN(n184) );
  AOI21_X1 U286 ( .B1(n563), .B2(n564), .A(n184), .ZN(n578) );
  NAND2_X1 U287 ( .A1(n186), .A2(n185), .ZN(n576) );
  FA_X1 U288 ( .A(n188), .B(f[4]), .CI(n187), .CO(n231), .S(n196) );
  XNOR2_X1 U289 ( .A(n664), .B(b_in[4]), .ZN(n190) );
  XNOR2_X1 U290 ( .A(b_in[5]), .B(a_in[0]), .ZN(n192) );
  INV_X1 U291 ( .A(n211), .ZN(n191) );
  XNOR2_X1 U292 ( .A(b_in[5]), .B(a_in[1]), .ZN(n213) );
  OAI22_X1 U293 ( .A1(n193), .A2(n192), .B1(n191), .B2(n213), .ZN(n216) );
  XNOR2_X1 U294 ( .A(n630), .B(a_in[5]), .ZN(n202) );
  OAI22_X1 U295 ( .A1(n299), .A2(n194), .B1(n202), .B2(n651), .ZN(n221) );
  XNOR2_X1 U296 ( .A(n633), .B(a_in[3]), .ZN(n215) );
  OAI22_X1 U297 ( .A1(n361), .A2(n195), .B1(n362), .B2(n215), .ZN(n220) );
  FA_X1 U298 ( .A(n198), .B(n197), .CI(n196), .CO(n199), .S(n186) );
  OR2_X1 U299 ( .A1(n200), .A2(n199), .ZN(n583) );
  NAND2_X1 U300 ( .A1(n200), .A2(n199), .ZN(n582) );
  INV_X1 U301 ( .A(n582), .ZN(n201) );
  XNOR2_X1 U302 ( .A(b_in[6]), .B(n664), .ZN(n206) );
  INV_X1 U303 ( .A(n206), .ZN(n208) );
  AND2_X1 U304 ( .A1(a_in[0]), .A2(n206), .ZN(n219) );
  XNOR2_X1 U305 ( .A(n630), .B(a_in[6]), .ZN(n203) );
  XNOR2_X1 U306 ( .A(n248), .B(a_in[7]), .ZN(n249) );
  OAI22_X1 U307 ( .A1(n299), .A2(n203), .B1(n249), .B2(n651), .ZN(n240) );
  XNOR2_X1 U308 ( .A(n431), .B(n639), .ZN(n205) );
  XNOR2_X1 U309 ( .A(n639), .B(n664), .ZN(n204) );
  XNOR2_X1 U310 ( .A(b_in[7]), .B(a_in[0]), .ZN(n207) );
  XNOR2_X1 U311 ( .A(b_in[7]), .B(a_in[1]), .ZN(n242) );
  OAI22_X1 U312 ( .A1(n140), .A2(n207), .B1(n435), .B2(n242), .ZN(n250) );
  INV_X1 U313 ( .A(b_in[7]), .ZN(n210) );
  OR2_X1 U314 ( .A1(a_in[0]), .A2(n210), .ZN(n209) );
  OAI22_X1 U315 ( .A1(n140), .A2(n210), .B1(n209), .B2(n435), .ZN(n253) );
  XNOR2_X1 U316 ( .A(b_in[5]), .B(a_in[2]), .ZN(n212) );
  XNOR2_X1 U317 ( .A(b_in[5]), .B(a_in[3]), .ZN(n247) );
  OAI22_X1 U318 ( .A1(n193), .A2(n212), .B1(n191), .B2(n247), .ZN(n252) );
  XNOR2_X1 U319 ( .A(n633), .B(a_in[4]), .ZN(n214) );
  XNOR2_X1 U320 ( .A(n633), .B(a_in[5]), .ZN(n246) );
  OAI22_X1 U321 ( .A1(n361), .A2(n214), .B1(n362), .B2(n246), .ZN(n251) );
  OAI22_X1 U322 ( .A1(n193), .A2(n213), .B1(n191), .B2(n212), .ZN(n225) );
  OAI22_X1 U323 ( .A1(n361), .A2(n215), .B1(n362), .B2(n214), .ZN(n224) );
  XNOR2_X1 U324 ( .A(n260), .B(n259), .ZN(n217) );
  FA_X1 U325 ( .A(n222), .B(n221), .CI(n220), .CO(n227), .S(n229) );
  FA_X1 U326 ( .A(n225), .B(n224), .CI(n223), .CO(n259), .S(n226) );
  FA_X1 U327 ( .A(n231), .B(n230), .CI(n229), .CO(n232), .S(n200) );
  NAND2_X1 U328 ( .A1(n597), .A2(n594), .ZN(n238) );
  INV_X1 U329 ( .A(n589), .ZN(n593) );
  INV_X1 U330 ( .A(n596), .ZN(n236) );
  OAI21_X1 U331 ( .B1(n588), .B2(n238), .A(n237), .ZN(n603) );
  FA_X1 U332 ( .A(n241), .B(n240), .CI(n239), .CO(n284), .S(n258) );
  INV_X1 U333 ( .A(n358), .ZN(n439) );
  XNOR2_X1 U334 ( .A(b_in[7]), .B(a_in[2]), .ZN(n267) );
  OR2_X1 U335 ( .A1(n435), .A2(n267), .ZN(n244) );
  NAND2_X1 U336 ( .A1(n245), .A2(n244), .ZN(n272) );
  XNOR2_X1 U337 ( .A(n633), .B(a_in[6]), .ZN(n279) );
  OAI22_X1 U338 ( .A1(n361), .A2(n246), .B1(n362), .B2(n279), .ZN(n271) );
  XNOR2_X1 U339 ( .A(b_in[5]), .B(a_in[4]), .ZN(n278) );
  OAI22_X1 U340 ( .A1(n193), .A2(n247), .B1(n359), .B2(n278), .ZN(n270) );
  XNOR2_X1 U341 ( .A(n663), .B(b_in[8]), .ZN(n264) );
  INV_X1 U342 ( .A(n264), .ZN(n321) );
  INV_X1 U343 ( .A(n321), .ZN(n386) );
  AND2_X1 U344 ( .A1(n386), .A2(a_in[0]), .ZN(n269) );
  XNOR2_X1 U345 ( .A(n248), .B(a_in[8]), .ZN(n266) );
  OAI22_X1 U346 ( .A1(n299), .A2(n249), .B1(n266), .B2(n651), .ZN(n268) );
  AND2_X1 U347 ( .A1(n250), .A2(f[7]), .ZN(n275) );
  XNOR2_X1 U348 ( .A(n274), .B(n275), .ZN(n254) );
  FA_X1 U349 ( .A(n252), .B(n251), .CI(n253), .CO(n273), .S(n260) );
  INV_X1 U350 ( .A(n260), .ZN(n256) );
  NAND2_X1 U351 ( .A1(n260), .A2(n259), .ZN(n261) );
  NOR2_X1 U352 ( .A1(n286), .A2(n285), .ZN(n602) );
  XNOR2_X1 U353 ( .A(n640), .B(n641), .ZN(n263) );
  OR2_X2 U354 ( .A1(n264), .A2(n263), .ZN(n445) );
  XNOR2_X1 U355 ( .A(n631), .B(a_in[0]), .ZN(n265) );
  XNOR2_X1 U356 ( .A(n631), .B(a_in[1]), .ZN(n294) );
  OAI22_X1 U357 ( .A1(n445), .A2(n265), .B1(n345), .B2(n294), .ZN(n306) );
  OAI22_X1 U358 ( .A1(n299), .A2(n266), .B1(n298), .B2(n651), .ZN(n305) );
  XNOR2_X1 U359 ( .A(b_in[7]), .B(a_in[3]), .ZN(n295) );
  OAI22_X1 U360 ( .A1(n358), .A2(n267), .B1(n208), .B2(n295), .ZN(n304) );
  FA_X1 U361 ( .A(n269), .B(f[8]), .CI(n268), .CO(n292), .S(n274) );
  FA_X1 U362 ( .A(n272), .B(n271), .CI(n270), .CO(n291), .S(n283) );
  OAI21_X1 U363 ( .B1(n275), .B2(n274), .A(n273), .ZN(n277) );
  NAND2_X1 U364 ( .A1(n277), .A2(n276), .ZN(n312) );
  XNOR2_X1 U365 ( .A(b_in[5]), .B(a_in[5]), .ZN(n302) );
  OAI22_X1 U366 ( .A1(n193), .A2(n278), .B1(n359), .B2(n302), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n633), .B(a_in[7]), .ZN(n325) );
  OAI22_X1 U368 ( .A1(n361), .A2(n279), .B1(n362), .B2(n325), .ZN(n308) );
  INV_X1 U369 ( .A(n631), .ZN(n280) );
  NAND2_X1 U370 ( .A1(n631), .A2(n144), .ZN(n281) );
  BUF_X1 U371 ( .A(n321), .Z(n345) );
  OAI22_X1 U372 ( .A1(n281), .A2(n345), .B1(n445), .B2(n280), .ZN(n296) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n282) );
  XNOR2_X1 U374 ( .A(n310), .B(n282), .ZN(n288) );
  NOR2_X1 U375 ( .A1(n288), .A2(n287), .ZN(n610) );
  NOR2_X1 U376 ( .A1(n602), .A2(n610), .ZN(n290) );
  NAND2_X1 U377 ( .A1(n288), .A2(n287), .ZN(n611) );
  INV_X1 U378 ( .A(n138), .ZN(n619) );
  XNOR2_X1 U379 ( .A(n136), .B(a_in[2]), .ZN(n322) );
  OAI22_X1 U380 ( .A1(n294), .A2(n445), .B1(n143), .B2(n322), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n431), .B(a_in[4]), .ZN(n318) );
  OAI22_X1 U382 ( .A1(n140), .A2(n295), .B1(n435), .B2(n318), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n633), .B(a_in[8]), .ZN(n324) );
  OAI22_X1 U384 ( .A1(n361), .A2(n325), .B1(n362), .B2(n324), .ZN(n301) );
  INV_X1 U385 ( .A(n300), .ZN(n327) );
  XNOR2_X1 U386 ( .A(n301), .B(n327), .ZN(n303) );
  XNOR2_X1 U387 ( .A(b_in[5]), .B(a_in[6]), .ZN(n319) );
  OAI22_X1 U388 ( .A1(n193), .A2(n302), .B1(n191), .B2(n319), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n303), .B(n328), .ZN(n317) );
  FA_X1 U390 ( .A(n305), .B(n306), .CI(n304), .CO(n316), .S(n293) );
  NAND2_X1 U391 ( .A1(n312), .A2(n311), .ZN(n313) );
  NAND2_X1 U392 ( .A1(n314), .A2(n313), .ZN(n406) );
  XNOR2_X1 U393 ( .A(b_in[7]), .B(a_in[5]), .ZN(n357) );
  OAI22_X1 U394 ( .A1(n140), .A2(n318), .B1(n435), .B2(n357), .ZN(n353) );
  XNOR2_X1 U395 ( .A(b_in[5]), .B(a_in[7]), .ZN(n360) );
  OAI22_X1 U396 ( .A1(n193), .A2(n319), .B1(n359), .B2(n360), .ZN(n352) );
  OR2_X1 U397 ( .A1(n320), .A2(f[10]), .ZN(n351) );
  XNOR2_X1 U398 ( .A(n136), .B(a_in[3]), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n348), .B(n145), .ZN(n323) );
  XNOR2_X1 U400 ( .A(n633), .B(a_in[9]), .ZN(n363) );
  OAI22_X1 U401 ( .A1(n362), .A2(n363), .B1(n361), .B2(n324), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n323), .B(n347), .ZN(n356) );
  OAI22_X1 U403 ( .A1(n361), .A2(n325), .B1(n362), .B2(n324), .ZN(n326) );
  OAI21_X1 U404 ( .B1(n328), .B2(n327), .A(n326), .ZN(n330) );
  OAI21_X1 U405 ( .B1(n333), .B2(n332), .A(n331), .ZN(n335) );
  NAND2_X1 U406 ( .A1(n335), .A2(n334), .ZN(n354) );
  OR2_X1 U407 ( .A1(n414), .A2(n413), .ZN(n379) );
  INV_X1 U408 ( .A(n379), .ZN(n344) );
  NAND2_X1 U409 ( .A1(n407), .A2(n406), .ZN(n341) );
  NAND2_X1 U410 ( .A1(n340), .A2(n339), .ZN(n408) );
  OAI21_X1 U411 ( .B1(n341), .B2(n342), .A(n408), .ZN(n425) );
  INV_X1 U412 ( .A(n425), .ZN(n376) );
  INV_X1 U413 ( .A(n376), .ZN(n343) );
  AOI21_X1 U414 ( .B1(n619), .B2(n344), .A(n343), .ZN(n374) );
  XNOR2_X1 U415 ( .A(n631), .B(a_in[4]), .ZN(n387) );
  OAI22_X1 U416 ( .A1(n445), .A2(n346), .B1(n345), .B2(n387), .ZN(n393) );
  OAI21_X1 U417 ( .B1(n142), .B2(n145), .A(n347), .ZN(n350) );
  NAND2_X1 U418 ( .A1(n142), .A2(n145), .ZN(n349) );
  FA_X1 U419 ( .A(n353), .B(n352), .CI(n351), .CO(n383), .S(n368) );
  FA_X1 U420 ( .A(n356), .B(n355), .CI(n354), .CO(n400), .S(n367) );
  XNOR2_X1 U421 ( .A(n431), .B(a_in[6]), .ZN(n392) );
  OAI22_X1 U422 ( .A1(n140), .A2(n357), .B1(n435), .B2(n392), .ZN(n391) );
  XNOR2_X1 U423 ( .A(b_in[5]), .B(a_in[8]), .ZN(n388) );
  OAI22_X1 U424 ( .A1(n193), .A2(n360), .B1(n359), .B2(n388), .ZN(n390) );
  NAND2_X1 U425 ( .A1(n362), .A2(n361), .ZN(n365) );
  INV_X1 U426 ( .A(n363), .ZN(n364) );
  NAND2_X1 U427 ( .A1(n365), .A2(n364), .ZN(n389) );
  XNOR2_X1 U428 ( .A(n400), .B(n399), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n398), .B(n366), .ZN(n371) );
  NOR2_X1 U430 ( .A1(n371), .A2(n370), .ZN(n418) );
  INV_X1 U431 ( .A(n378), .ZN(n372) );
  NAND2_X1 U432 ( .A1(n371), .A2(n370), .ZN(n421) );
  INV_X1 U433 ( .A(reset), .ZN(n540) );
  NOR2_X2 U434 ( .A1(enable_f), .A2(reset), .ZN(n627) );
  NAND2_X1 U435 ( .A1(n627), .A2(f[12]), .ZN(n375) );
  OAI21_X1 U436 ( .B1(n376), .B2(n378), .A(n421), .ZN(n377) );
  INV_X1 U437 ( .A(n377), .ZN(n382) );
  NOR2_X1 U438 ( .A1(n379), .A2(n378), .ZN(n380) );
  NAND2_X1 U439 ( .A1(n619), .A2(n380), .ZN(n381) );
  FA_X1 U440 ( .A(n385), .B(n384), .CI(n383), .CO(n471), .S(n398) );
  XNOR2_X1 U441 ( .A(n631), .B(a_in[5]), .ZN(n444) );
  OAI22_X1 U442 ( .A1(n445), .A2(n387), .B1(n426), .B2(n444), .ZN(n452) );
  XNOR2_X1 U443 ( .A(b_in[5]), .B(a_in[9]), .ZN(n446) );
  OAI22_X1 U444 ( .A1(n193), .A2(n388), .B1(n359), .B2(n446), .ZN(n451) );
  FA_X1 U445 ( .A(n391), .B(n390), .CI(n389), .CO(n464), .S(n399) );
  INV_X1 U446 ( .A(n439), .ZN(n450) );
  XNOR2_X1 U447 ( .A(b_in[7]), .B(a_in[7]), .ZN(n449) );
  FA_X1 U448 ( .A(f[11]), .B(f[12]), .CI(n393), .CO(n465), .S(n385) );
  XNOR2_X1 U449 ( .A(n466), .B(n465), .ZN(n394) );
  INV_X1 U450 ( .A(n400), .ZN(n396) );
  INV_X1 U451 ( .A(n399), .ZN(n395) );
  NAND2_X1 U452 ( .A1(n396), .A2(n395), .ZN(n397) );
  NAND2_X1 U453 ( .A1(n398), .A2(n397), .ZN(n402) );
  NAND2_X1 U454 ( .A1(n402), .A2(n401), .ZN(n415) );
  NOR2_X1 U455 ( .A1(n416), .A2(n415), .ZN(n422) );
  INV_X1 U456 ( .A(n417), .ZN(n403) );
  NAND2_X1 U457 ( .A1(n416), .A2(n415), .ZN(n420) );
  NAND2_X1 U458 ( .A1(n627), .A2(f[13]), .ZN(n404) );
  OAI21_X1 U459 ( .B1(n405), .B2(n499), .A(n404), .ZN(n54) );
  AND2_X1 U460 ( .A1(n407), .A2(n406), .ZN(n616) );
  AOI21_X1 U461 ( .B1(n619), .B2(n137), .A(n616), .ZN(n410) );
  NAND2_X1 U462 ( .A1(n141), .A2(n408), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n410), .B(n409), .ZN(n412) );
  NOR2_X1 U464 ( .A1(n416), .A2(n415), .ZN(n417) );
  NOR2_X1 U465 ( .A1(n418), .A2(n417), .ZN(n424) );
  NAND2_X1 U466 ( .A1(n419), .A2(n424), .ZN(n510) );
  OAI21_X1 U467 ( .B1(n422), .B2(n421), .A(n420), .ZN(n423) );
  AOI21_X1 U468 ( .B1(n425), .B2(n424), .A(n423), .ZN(n509) );
  OAI21_X1 U469 ( .B1(n138), .B2(n510), .A(n509), .ZN(n626) );
  XNOR2_X1 U470 ( .A(n631), .B(a_in[8]), .ZN(n427) );
  XNOR2_X1 U471 ( .A(n631), .B(a_in[9]), .ZN(n428) );
  OAI22_X1 U472 ( .A1(n445), .A2(n427), .B1(n426), .B2(n428), .ZN(n454) );
  XNOR2_X1 U473 ( .A(n631), .B(a_in[7]), .ZN(n430) );
  OAI22_X1 U474 ( .A1(n445), .A2(n430), .B1(n426), .B2(n427), .ZN(n440) );
  AOI21_X1 U475 ( .B1(n426), .B2(n445), .A(n428), .ZN(n429) );
  INV_X1 U476 ( .A(n429), .ZN(n479) );
  OR2_X1 U477 ( .A1(n496), .A2(n495), .ZN(n516) );
  XNOR2_X1 U478 ( .A(n631), .B(a_in[6]), .ZN(n443) );
  OAI22_X1 U479 ( .A1(n443), .A2(n445), .B1(n426), .B2(n430), .ZN(n442) );
  XNOR2_X1 U480 ( .A(n431), .B(a_in[8]), .ZN(n448) );
  INV_X1 U481 ( .A(n448), .ZN(n432) );
  NAND2_X1 U482 ( .A1(n439), .A2(n432), .ZN(n434) );
  XNOR2_X1 U483 ( .A(b_in[7]), .B(a_in[9]), .ZN(n436) );
  OR2_X1 U484 ( .A1(n435), .A2(n436), .ZN(n433) );
  NAND2_X1 U485 ( .A1(n434), .A2(n433), .ZN(n441) );
  INV_X1 U486 ( .A(n435), .ZN(n438) );
  INV_X1 U487 ( .A(n436), .ZN(n437) );
  OAI21_X1 U488 ( .B1(n439), .B2(n438), .A(n437), .ZN(n456) );
  FA_X1 U489 ( .A(f[15]), .B(f[16]), .CI(n440), .CO(n453), .S(n455) );
  FA_X1 U490 ( .A(n442), .B(n650), .CI(n441), .CO(n457), .S(n474) );
  OAI22_X1 U491 ( .A1(n445), .A2(n444), .B1(n426), .B2(n443), .ZN(n462) );
  AOI21_X1 U492 ( .B1(n193), .B2(n359), .A(n446), .ZN(n447) );
  INV_X1 U493 ( .A(n447), .ZN(n461) );
  OAI22_X1 U494 ( .A1(n450), .A2(n449), .B1(n435), .B2(n448), .ZN(n460) );
  FA_X1 U495 ( .A(n452), .B(n146), .CI(n451), .CO(n459), .S(n470) );
  NOR2_X1 U496 ( .A1(n489), .A2(n488), .ZN(n526) );
  INV_X1 U497 ( .A(n526), .ZN(n521) );
  FA_X1 U498 ( .A(n454), .B(n649), .CI(n453), .CO(n496), .S(n491) );
  FA_X1 U499 ( .A(n457), .B(n456), .CI(n455), .CO(n490), .S(n489) );
  OR2_X1 U500 ( .A1(n491), .A2(n490), .ZN(n531) );
  NAND2_X1 U501 ( .A1(n521), .A2(n531), .ZN(n512) );
  INV_X1 U502 ( .A(n512), .ZN(n458) );
  NAND2_X1 U503 ( .A1(n516), .A2(n458), .ZN(n478) );
  FA_X1 U504 ( .A(f[13]), .B(f[14]), .CI(n462), .CO(n473), .S(n476) );
  OR2_X1 U505 ( .A1(n465), .A2(n466), .ZN(n463) );
  NAND2_X1 U506 ( .A1(n466), .A2(n465), .ZN(n467) );
  OR2_X1 U507 ( .A1(n484), .A2(n483), .ZN(n624) );
  FA_X1 U508 ( .A(n474), .B(n473), .CI(n472), .CO(n488), .S(n486) );
  FA_X1 U509 ( .A(n477), .B(n476), .CI(n475), .CO(n485), .S(n484) );
  OR2_X1 U510 ( .A1(n486), .A2(n485), .ZN(n536) );
  NAND2_X1 U511 ( .A1(n624), .A2(n536), .ZN(n524) );
  NOR2_X1 U512 ( .A1(n478), .A2(n524), .ZN(n502) );
  FA_X1 U513 ( .A(f[17]), .B(f[18]), .CI(n479), .CO(n480), .S(n495) );
  OR2_X1 U514 ( .A1(n480), .A2(n648), .ZN(n482) );
  NAND2_X1 U515 ( .A1(n480), .A2(n648), .ZN(n481) );
  AND2_X1 U516 ( .A1(n482), .A2(n481), .ZN(n503) );
  NAND2_X1 U517 ( .A1(n626), .A2(n152), .ZN(n501) );
  AND2_X2 U518 ( .A1(n484), .A2(n483), .ZN(n622) );
  NAND2_X1 U519 ( .A1(n486), .A2(n485), .ZN(n535) );
  INV_X1 U520 ( .A(n535), .ZN(n487) );
  NAND2_X1 U521 ( .A1(n489), .A2(n488), .ZN(n525) );
  INV_X1 U522 ( .A(n525), .ZN(n493) );
  NAND2_X1 U523 ( .A1(n491), .A2(n490), .ZN(n530) );
  INV_X1 U524 ( .A(n530), .ZN(n492) );
  AOI21_X1 U525 ( .B1(n493), .B2(n531), .A(n492), .ZN(n494) );
  OAI21_X1 U526 ( .B1(n527), .B2(n512), .A(n494), .ZN(n513) );
  NAND2_X1 U527 ( .A1(n496), .A2(n495), .ZN(n515) );
  INV_X1 U528 ( .A(n515), .ZN(n497) );
  AOI21_X1 U529 ( .B1(n513), .B2(n516), .A(n497), .ZN(n498) );
  INV_X1 U530 ( .A(n665), .ZN(n499) );
  AOI21_X1 U531 ( .B1(n626), .B2(n502), .A(n503), .ZN(n507) );
  NAND2_X1 U532 ( .A1(n627), .A2(f[19]), .ZN(n506) );
  INV_X1 U533 ( .A(n503), .ZN(n504) );
  NAND2_X1 U534 ( .A1(n504), .A2(n665), .ZN(n505) );
  OAI211_X1 U535 ( .C1(n508), .C2(n507), .A(n506), .B(n158), .ZN(n48) );
  OAI21_X1 U536 ( .B1(n510), .B2(n511), .A(n509), .ZN(n534) );
  NOR2_X1 U537 ( .A1(n524), .A2(n512), .ZN(n514) );
  AOI21_X1 U538 ( .B1(n534), .B2(n514), .A(n513), .ZN(n517) );
  XNOR2_X1 U539 ( .A(n517), .B(n149), .ZN(n518) );
  OAI21_X1 U540 ( .B1(n518), .B2(n499), .A(n154), .ZN(n49) );
  INV_X1 U541 ( .A(n524), .ZN(n520) );
  INV_X1 U542 ( .A(n527), .ZN(n519) );
  AOI21_X1 U543 ( .B1(n534), .B2(n520), .A(n519), .ZN(n522) );
  XNOR2_X1 U544 ( .A(n522), .B(n148), .ZN(n523) );
  OAI21_X1 U545 ( .B1(n523), .B2(n499), .A(n155), .ZN(n51) );
  NOR2_X1 U546 ( .A1(n524), .A2(n526), .ZN(n529) );
  OAI21_X1 U547 ( .B1(n527), .B2(n526), .A(n525), .ZN(n528) );
  AOI21_X1 U548 ( .B1(n534), .B2(n529), .A(n528), .ZN(n532) );
  XNOR2_X1 U549 ( .A(n532), .B(n150), .ZN(n533) );
  OAI21_X1 U550 ( .B1(n533), .B2(n499), .A(n156), .ZN(n50) );
  AOI21_X1 U551 ( .B1(n534), .B2(n624), .A(n622), .ZN(n537) );
  XNOR2_X1 U552 ( .A(n537), .B(n151), .ZN(n538) );
  OAI21_X1 U553 ( .B1(n538), .B2(n499), .A(n157), .ZN(n52) );
  INV_X1 U554 ( .A(n635), .ZN(n539) );
  OAI21_X1 U555 ( .B1(n652), .B2(n540), .A(n539), .ZN(n47) );
  OR2_X1 U556 ( .A1(n541), .A2(f[0]), .ZN(n542) );
  AND2_X1 U557 ( .A1(n542), .A2(n558), .ZN(n543) );
  AOI22_X1 U558 ( .A1(n543), .A2(n665), .B1(n627), .B2(f[0]), .ZN(n544) );
  INV_X1 U559 ( .A(n544), .ZN(n67) );
  NOR2_X2 U560 ( .A1(valid_in), .A2(reset), .ZN(n634) );
  AOI22_X1 U561 ( .A1(n635), .A2(a[9]), .B1(n634), .B2(a_in[9]), .ZN(n545) );
  INV_X1 U562 ( .A(n545), .ZN(n77) );
  AOI22_X1 U563 ( .A1(n635), .A2(a[7]), .B1(n634), .B2(a_in[7]), .ZN(n546) );
  INV_X1 U564 ( .A(n546), .ZN(n79) );
  AOI22_X1 U565 ( .A1(n635), .A2(a[8]), .B1(n634), .B2(a_in[8]), .ZN(n547) );
  INV_X1 U566 ( .A(n547), .ZN(n78) );
  AOI22_X1 U567 ( .A1(n635), .A2(a[6]), .B1(n634), .B2(a_in[6]), .ZN(n548) );
  INV_X1 U568 ( .A(n548), .ZN(n80) );
  AOI22_X1 U569 ( .A1(n635), .A2(a[5]), .B1(n634), .B2(a_in[5]), .ZN(n549) );
  INV_X1 U570 ( .A(n549), .ZN(n81) );
  AOI22_X1 U571 ( .A1(n635), .A2(a[4]), .B1(n634), .B2(a_in[4]), .ZN(n656) );
  AOI22_X1 U572 ( .A1(n635), .A2(a[3]), .B1(n634), .B2(a_in[3]), .ZN(n550) );
  INV_X1 U573 ( .A(n550), .ZN(n83) );
  AOI22_X1 U574 ( .A1(n635), .A2(b[8]), .B1(n634), .B2(b_in[8]), .ZN(n657) );
  AOI22_X1 U575 ( .A1(n635), .A2(a[2]), .B1(n634), .B2(a_in[2]), .ZN(n551) );
  INV_X1 U576 ( .A(n551), .ZN(n84) );
  AOI22_X1 U577 ( .A1(n635), .A2(a[1]), .B1(n634), .B2(a_in[1]), .ZN(n552) );
  INV_X1 U578 ( .A(n552), .ZN(n85) );
  AOI22_X1 U579 ( .A1(n635), .A2(a[0]), .B1(n634), .B2(a_in[0]), .ZN(n553) );
  INV_X1 U580 ( .A(n553), .ZN(n86) );
  AOI22_X1 U581 ( .A1(n635), .A2(b[6]), .B1(n634), .B2(b_in[6]), .ZN(n658) );
  AOI22_X1 U582 ( .A1(n635), .A2(b[4]), .B1(n634), .B2(b_in[4]), .ZN(n554) );
  INV_X1 U583 ( .A(n554), .ZN(n73) );
  AOI22_X1 U584 ( .A1(n635), .A2(b[2]), .B1(n634), .B2(b_in[2]), .ZN(n659) );
  AOI22_X1 U585 ( .A1(n635), .A2(b[0]), .B1(n634), .B2(b_in[0]), .ZN(n660) );
  INV_X1 U586 ( .A(n555), .ZN(n557) );
  NAND2_X1 U587 ( .A1(n557), .A2(n556), .ZN(n559) );
  XOR2_X1 U588 ( .A(n559), .B(n558), .Z(n560) );
  AOI22_X1 U589 ( .A1(n560), .A2(n665), .B1(n627), .B2(f[1]), .ZN(n561) );
  INV_X1 U590 ( .A(n561), .ZN(n66) );
  NAND2_X1 U591 ( .A1(n563), .A2(n562), .ZN(n565) );
  XNOR2_X1 U592 ( .A(n565), .B(n564), .ZN(n566) );
  AOI22_X1 U593 ( .A1(n566), .A2(n665), .B1(n627), .B2(f[3]), .ZN(n567) );
  INV_X1 U594 ( .A(n567), .ZN(n64) );
  INV_X1 U595 ( .A(n568), .ZN(n570) );
  NAND2_X1 U596 ( .A1(n570), .A2(n569), .ZN(n572) );
  XOR2_X1 U597 ( .A(n572), .B(n571), .Z(n573) );
  AOI22_X1 U598 ( .A1(n573), .A2(n665), .B1(n627), .B2(f[2]), .ZN(n574) );
  INV_X1 U599 ( .A(n574), .ZN(n65) );
  INV_X1 U600 ( .A(n575), .ZN(n577) );
  NAND2_X1 U601 ( .A1(n577), .A2(n576), .ZN(n579) );
  XOR2_X1 U602 ( .A(n578), .B(n579), .Z(n580) );
  AOI22_X1 U603 ( .A1(n580), .A2(n665), .B1(n627), .B2(f[4]), .ZN(n581) );
  INV_X1 U604 ( .A(n581), .ZN(n63) );
  NAND2_X1 U605 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U606 ( .A(n585), .B(n584), .ZN(n586) );
  AOI22_X1 U607 ( .A1(n586), .A2(n665), .B1(n627), .B2(f[5]), .ZN(n587) );
  INV_X1 U608 ( .A(n587), .ZN(n62) );
  INV_X1 U609 ( .A(n588), .ZN(n595) );
  NAND2_X1 U610 ( .A1(n594), .A2(n589), .ZN(n590) );
  XNOR2_X1 U611 ( .A(n595), .B(n590), .ZN(n591) );
  AOI22_X1 U612 ( .A1(n591), .A2(n665), .B1(n627), .B2(f[6]), .ZN(n592) );
  INV_X1 U613 ( .A(n592), .ZN(n61) );
  AOI21_X1 U614 ( .B1(n595), .B2(n594), .A(n593), .ZN(n599) );
  NAND2_X1 U615 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U616 ( .A(n599), .B(n598), .Z(n600) );
  AOI22_X1 U617 ( .A1(n600), .A2(n665), .B1(n627), .B2(f[7]), .ZN(n601) );
  INV_X1 U618 ( .A(n601), .ZN(n60) );
  INV_X1 U619 ( .A(n602), .ZN(n606) );
  NAND2_X1 U620 ( .A1(n606), .A2(n607), .ZN(n604) );
  INV_X1 U621 ( .A(n139), .ZN(n609) );
  XOR2_X1 U622 ( .A(n604), .B(n609), .Z(n605) );
  AOI22_X1 U623 ( .A1(n605), .A2(n665), .B1(n627), .B2(f[8]), .ZN(n662) );
  INV_X1 U624 ( .A(n606), .ZN(n608) );
  OAI21_X1 U625 ( .B1(n609), .B2(n608), .A(n607), .ZN(n614) );
  INV_X1 U626 ( .A(n610), .ZN(n612) );
  NAND2_X1 U627 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U628 ( .A(n614), .B(n613), .ZN(n615) );
  AOI22_X1 U629 ( .A1(n615), .A2(n665), .B1(n627), .B2(f[9]), .ZN(n661) );
  INV_X1 U630 ( .A(n616), .ZN(n617) );
  NAND2_X1 U631 ( .A1(n137), .A2(n617), .ZN(n618) );
  XNOR2_X1 U632 ( .A(n619), .B(n618), .ZN(n620) );
  AOI22_X1 U633 ( .A1(n620), .A2(n665), .B1(n627), .B2(f[10]), .ZN(n621) );
  INV_X1 U634 ( .A(n621), .ZN(n57) );
  INV_X1 U635 ( .A(n622), .ZN(n623) );
  NAND2_X1 U636 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U637 ( .A(n626), .B(n625), .ZN(n628) );
  AOI22_X1 U638 ( .A1(n628), .A2(n665), .B1(n627), .B2(f[14]), .ZN(n629) );
  INV_X1 U639 ( .A(n629), .ZN(n53) );
  AOI22_X1 U640 ( .A1(n635), .A2(b[1]), .B1(n634), .B2(n630), .ZN(n653) );
  AOI22_X1 U641 ( .A1(n635), .A2(b[9]), .B1(n634), .B2(n631), .ZN(n654) );
  AOI22_X1 U642 ( .A1(n635), .A2(b[5]), .B1(n634), .B2(b_in[5]), .ZN(n632) );
  INV_X1 U643 ( .A(n632), .ZN(n72) );
  AOI22_X1 U644 ( .A1(n635), .A2(b[3]), .B1(n634), .B2(n633), .ZN(n655) );
  AOI22_X1 U645 ( .A1(n635), .A2(b[7]), .B1(n634), .B2(b_in[7]), .ZN(n636) );
  INV_X1 U646 ( .A(n636), .ZN(n70) );
endmodule

