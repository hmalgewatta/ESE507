
module part1_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   enable_f, n45, n46, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n68, n70, n73, n84,
         \DP_OP_12J1_122_830/n469 , n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789;
  wire   [9:0] a_in;
  wire   [9:0] b_in;

  DFF_X1 enable_f_reg ( .D(n134), .CK(clk), .Q(enable_f), .QN(n773) );
  DFF_X1 \f_reg[17]  ( .D(n47), .CK(clk), .Q(f[17]) );
  DFF_X1 \f_reg[16]  ( .D(n48), .CK(clk), .Q(f[16]), .QN(n138) );
  DFF_X1 \f_reg[14]  ( .D(n50), .CK(clk), .Q(f[14]), .QN(n136) );
  DFF_X1 \f_reg[13]  ( .D(n51), .CK(clk), .Q(f[13]) );
  DFF_X1 \f_reg[12]  ( .D(n52), .CK(clk), .Q(f[12]) );
  DFF_X1 \f_reg[11]  ( .D(n53), .CK(clk), .Q(f[11]) );
  DFF_X1 \b_in_reg[9]  ( .D(n65), .CK(clk), .Q(b_in[9]), .QN(n142) );
  DFF_X1 \b_in_reg[8]  ( .D(n66), .CK(clk), .Q(b_in[8]), .QN(n141) );
  DFF_X1 \b_in_reg[4]  ( .D(n70), .CK(clk), .Q(b_in[4]), .QN(n140) );
  DFF_X1 \b_in_reg[1]  ( .D(n73), .CK(clk), .Q(b_in[1]), .QN(n139) );
  DFF_X1 \f_reg[19]  ( .D(n45), .CK(clk), .Q(f[19]) );
  DFF_X1 \a_in_reg[3]  ( .D(n775), .CK(clk), .Q(n760), .QN(
        \DP_OP_12J1_122_830/n469 ) );
  DFF_X1 \a_in_reg[5]  ( .D(n776), .CK(clk), .Q(n759), .QN(a_in[5]) );
  DFF_X1 \a_in_reg[1]  ( .D(n778), .CK(clk), .Q(n762), .QN(a_in[1]) );
  DFF_X1 \a_in_reg[2]  ( .D(n782), .CK(clk), .Q(n771), .QN(a_in[2]) );
  DFF_X1 \a_in_reg[7]  ( .D(n777), .CK(clk), .Q(n758), .QN(a_in[7]) );
  DFF_X1 \a_in_reg[4]  ( .D(n781), .CK(clk), .Q(n772), .QN(a_in[4]) );
  DFF_X1 valid_out_reg ( .D(n789), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[0]  ( .D(n64), .CK(clk), .Q(f[0]) );
  DFF_X1 \b_in_reg[6]  ( .D(n68), .CK(clk), .Q(b_in[6]), .QN(n767) );
  DFF_X1 \f_reg[1]  ( .D(n63), .CK(clk), .Q(f[1]) );
  DFF_X1 \f_reg[2]  ( .D(n62), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(n61), .CK(clk), .Q(f[3]) );
  DFF_X1 \f_reg[4]  ( .D(n60), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(n59), .CK(clk), .Q(f[5]) );
  DFF_X1 \f_reg[6]  ( .D(n58), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(n57), .CK(clk), .Q(f[7]), .QN(n756) );
  DFF_X1 \f_reg[8]  ( .D(n56), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[9]  ( .D(n55), .CK(clk), .Q(f[9]), .QN(n763) );
  DFF_X1 \a_in_reg[6]  ( .D(n780), .CK(clk), .QN(a_in[6]) );
  DFF_X1 \f_reg[10]  ( .D(n788), .CK(clk), .QN(f[10]) );
  DFF_X1 \a_in_reg[0]  ( .D(n783), .CK(clk), .Q(n769), .QN(a_in[0]) );
  DFF_X1 \b_in_reg[3]  ( .D(n786), .CK(clk), .Q(n770), .QN(b_in[3]) );
  DFF_X1 \b_in_reg[5]  ( .D(n785), .CK(clk), .Q(n768), .QN(b_in[5]) );
  DFF_X1 \b_in_reg[7]  ( .D(n784), .CK(clk), .Q(n766), .QN(b_in[7]) );
  SDFF_X1 \a_in_reg[8]  ( .D(n779), .SI(1'b0), .SE(1'b0), .CK(clk), .Q(n757), 
        .QN(a_in[8]) );
  SDFFRS_X2 \b_in_reg[2]  ( .D(n787), .SI(1'b0), .SE(1'b0), .CK(clk), .RN(1'b1), .SN(1'b1), .QN(b_in[2]) );
  DFF_X1 \a_in_reg[9]  ( .D(n774), .CK(clk), .Q(n764), .QN(a_in[9]) );
  DFF_X1 \b_in_reg[0]  ( .D(n84), .CK(clk), .Q(b_in[0]), .QN(n761) );
  DFF_X1 \f_reg[18]  ( .D(n46), .CK(clk), .Q(f[18]), .QN(n765) );
  DFF_X1 \f_reg[15]  ( .D(n49), .CK(clk), .Q(f[15]) );
  BUF_X1 U89 ( .A(a_in[5]), .Z(n114) );
  OAI22_X1 U90 ( .A1(n133), .A2(n196), .B1(n420), .B2(n163), .ZN(n228) );
  OAI21_X1 U91 ( .B1(n603), .B2(n606), .A(n604), .ZN(n623) );
  AND2_X2 U92 ( .A1(n288), .A2(n287), .ZN(n701) );
  CLKBUF_X1 U93 ( .A(n671), .Z(n672) );
  OR2_X1 U94 ( .A1(n529), .A2(n528), .ZN(n120) );
  AND2_X1 U95 ( .A1(n319), .A2(n318), .ZN(n95) );
  BUF_X1 U96 ( .A(b_in[2]), .Z(n111) );
  NAND2_X1 U97 ( .A1(n477), .A2(n476), .ZN(n478) );
  INV_X1 U98 ( .A(n480), .ZN(n476) );
  INV_X1 U99 ( .A(n389), .ZN(n385) );
  INV_X1 U100 ( .A(n388), .ZN(n384) );
  OR2_X1 U101 ( .A1(n434), .A2(f[13]), .ZN(n432) );
  NAND2_X1 U102 ( .A1(n434), .A2(f[13]), .ZN(n435) );
  NAND2_X1 U103 ( .A1(n496), .A2(n495), .ZN(n497) );
  NAND2_X1 U104 ( .A1(n494), .A2(n493), .ZN(n495) );
  OAI21_X1 U105 ( .B1(n494), .B2(n493), .A(n492), .ZN(n496) );
  NAND2_X1 U106 ( .A1(n437), .A2(n136), .ZN(n425) );
  OR2_X1 U107 ( .A1(n437), .A2(n136), .ZN(n424) );
  NAND2_X1 U108 ( .A1(n286), .A2(n285), .ZN(n407) );
  NAND2_X1 U109 ( .A1(n399), .A2(n143), .ZN(n286) );
  CLKBUF_X1 U110 ( .A(n644), .Z(n630) );
  CLKBUF_X1 U111 ( .A(n693), .Z(n118) );
  NAND2_X1 U112 ( .A1(n531), .A2(n789), .ZN(n541) );
  INV_X1 U113 ( .A(n536), .ZN(n531) );
  AND2_X1 U114 ( .A1(n537), .A2(n146), .ZN(n538) );
  CLKBUF_X1 U115 ( .A(a_in[5]), .Z(n750) );
  CLKBUF_X1 U116 ( .A(n189), .Z(n124) );
  CLKBUF_X1 U117 ( .A(n380), .Z(n125) );
  CLKBUF_X1 U118 ( .A(n759), .Z(n126) );
  NAND2_X1 U119 ( .A1(n352), .A2(n351), .ZN(n353) );
  NAND2_X1 U120 ( .A1(n348), .A2(n347), .ZN(n352) );
  BUF_X1 U121 ( .A(a_in[1]), .Z(n335) );
  CLKBUF_X1 U122 ( .A(n484), .Z(n525) );
  CLKBUF_X1 U123 ( .A(n244), .Z(n87) );
  XNOR2_X1 U124 ( .A(n243), .B(n242), .ZN(n245) );
  CLKBUF_X1 U125 ( .A(n246), .Z(n250) );
  NAND2_X1 U126 ( .A1(n441), .A2(n440), .ZN(n442) );
  XNOR2_X1 U127 ( .A(n437), .B(n136), .ZN(n438) );
  INV_X1 U128 ( .A(n262), .ZN(n258) );
  NAND2_X1 U129 ( .A1(n389), .A2(n388), .ZN(n390) );
  NAND2_X1 U130 ( .A1(n385), .A2(n384), .ZN(n387) );
  AND2_X1 U131 ( .A1(n354), .A2(n353), .ZN(n643) );
  XNOR2_X1 U132 ( .A(n348), .B(n294), .ZN(n334) );
  CLKBUF_X1 U133 ( .A(n760), .Z(n104) );
  NAND2_X1 U134 ( .A1(n436), .A2(n435), .ZN(n461) );
  XNOR2_X1 U135 ( .A(n434), .B(f[13]), .ZN(n154) );
  NAND2_X1 U136 ( .A1(n483), .A2(n482), .ZN(n517) );
  NAND2_X1 U137 ( .A1(n481), .A2(n480), .ZN(n482) );
  CLKBUF_X1 U138 ( .A(n655), .Z(n656) );
  CLKBUF_X1 U139 ( .A(n737), .Z(n567) );
  INV_X1 U140 ( .A(n568), .ZN(n560) );
  CLKBUF_X1 U141 ( .A(n670), .Z(n109) );
  CLKBUF_X1 U142 ( .A(n665), .Z(n107) );
  CLKBUF_X1 U143 ( .A(n657), .Z(n662) );
  CLKBUF_X1 U144 ( .A(n653), .Z(n654) );
  CLKBUF_X1 U145 ( .A(n616), .Z(n130) );
  CLKBUF_X1 U146 ( .A(n620), .Z(n97) );
  INV_X1 U147 ( .A(n95), .ZN(n610) );
  CLKBUF_X1 U148 ( .A(n513), .Z(n129) );
  AND2_X1 U149 ( .A1(n503), .A2(n789), .ZN(n504) );
  CLKBUF_X1 U150 ( .A(n645), .Z(n632) );
  CLKBUF_X1 U151 ( .A(n635), .Z(n640) );
  CLKBUF_X1 U152 ( .A(a_in[4]), .Z(n112) );
  NAND2_X1 U153 ( .A1(n688), .A2(n789), .ZN(n690) );
  NAND2_X1 U154 ( .A1(n696), .A2(n789), .ZN(n698) );
  OAI21_X1 U155 ( .B1(n537), .B2(n541), .A(n534), .ZN(n535) );
  NAND2_X1 U156 ( .A1(n178), .A2(n177), .ZN(n85) );
  XNOR2_X1 U157 ( .A(n758), .B(n757), .ZN(n86) );
  INV_X1 U158 ( .A(n102), .ZN(n751) );
  OR2_X1 U159 ( .A1(n401), .A2(n404), .ZN(n88) );
  OR2_X1 U160 ( .A1(n502), .A2(n706), .ZN(n89) );
  XNOR2_X1 U161 ( .A(n256), .B(n255), .ZN(n90) );
  INV_X1 U162 ( .A(n141), .ZN(n91) );
  BUF_X2 U163 ( .A(a_in[1]), .Z(n92) );
  XNOR2_X1 U164 ( .A(n386), .B(n367), .ZN(n372) );
  XNOR2_X1 U165 ( .A(n324), .B(n323), .ZN(n326) );
  XNOR2_X1 U166 ( .A(n326), .B(n325), .ZN(n331) );
  INV_X1 U167 ( .A(n535), .ZN(n540) );
  NOR2_X2 U168 ( .A1(n475), .A2(n474), .ZN(n706) );
  NAND2_X1 U169 ( .A1(n281), .A2(n280), .ZN(n93) );
  INV_X1 U170 ( .A(n629), .ZN(n94) );
  INV_X1 U171 ( .A(n643), .ZN(n629) );
  XOR2_X1 U172 ( .A(n762), .B(b_in[7]), .Z(n356) );
  INV_X1 U173 ( .A(n760), .ZN(n96) );
  BUF_X2 U174 ( .A(\DP_OP_12J1_122_830/n469 ), .Z(n749) );
  OAI21_X1 U175 ( .B1(n444), .B2(n443), .A(n442), .ZN(n464) );
  NOR2_X1 U176 ( .A1(n441), .A2(n440), .ZN(n444) );
  OAI21_X1 U177 ( .B1(n122), .B2(n159), .A(n158), .ZN(n441) );
  XOR2_X1 U178 ( .A(n228), .B(n227), .Z(n98) );
  XOR2_X1 U179 ( .A(n229), .B(n98), .Z(n262) );
  NAND2_X1 U180 ( .A1(n229), .A2(n228), .ZN(n99) );
  NAND2_X1 U181 ( .A1(n229), .A2(n227), .ZN(n100) );
  NAND2_X1 U182 ( .A1(n228), .A2(n227), .ZN(n101) );
  NAND3_X1 U183 ( .A1(n99), .A2(n100), .A3(n101), .ZN(n185) );
  INV_X1 U184 ( .A(n762), .ZN(n102) );
  XNOR2_X1 U185 ( .A(n245), .B(n87), .ZN(n264) );
  NAND2_X1 U186 ( .A1(n205), .A2(n155), .ZN(n103) );
  OAI21_X1 U187 ( .B1(n706), .B2(n702), .A(n707), .ZN(n105) );
  INV_X1 U188 ( .A(n309), .ZN(n342) );
  INV_X1 U189 ( .A(n213), .ZN(n106) );
  OR2_X1 U190 ( .A1(n354), .A2(n353), .ZN(n644) );
  NAND2_X1 U191 ( .A1(n281), .A2(n280), .ZN(n393) );
  INV_X1 U192 ( .A(n761), .ZN(n108) );
  NOR2_X1 U193 ( .A1(n415), .A2(n414), .ZN(n110) );
  XOR2_X1 U194 ( .A(n102), .B(n768), .Z(n336) );
  OR2_X2 U195 ( .A1(n174), .A2(n309), .ZN(n113) );
  OR2_X1 U196 ( .A1(n174), .A2(n309), .ZN(n344) );
  NOR2_X1 U197 ( .A1(n408), .A2(n407), .ZN(n670) );
  BUF_X2 U198 ( .A(a_in[5]), .Z(n115) );
  NAND2_X1 U199 ( .A1(n412), .A2(n411), .ZN(n116) );
  NAND3_X1 U200 ( .A1(n511), .A2(n506), .A3(n504), .ZN(n509) );
  BUF_X1 U201 ( .A(n309), .Z(n117) );
  NOR2_X1 U202 ( .A1(n529), .A2(n528), .ZN(n119) );
  NOR2_X1 U203 ( .A1(n529), .A2(n528), .ZN(n562) );
  XNOR2_X1 U204 ( .A(n233), .B(n260), .ZN(n121) );
  BUF_X1 U205 ( .A(n204), .Z(n122) );
  BUF_X1 U206 ( .A(n204), .Z(n722) );
  NAND2_X1 U207 ( .A1(n216), .A2(n215), .ZN(n123) );
  NOR2_X1 U208 ( .A1(n205), .A2(n761), .ZN(n275) );
  AND2_X1 U209 ( .A1(n224), .A2(f[9]), .ZN(n243) );
  INV_X1 U210 ( .A(n721), .ZN(n127) );
  INV_X1 U211 ( .A(n127), .ZN(n128) );
  BUF_X2 U212 ( .A(n149), .Z(n524) );
  NAND2_X1 U213 ( .A1(n350), .A2(n349), .ZN(n351) );
  OR2_X1 U214 ( .A1(n350), .A2(n349), .ZN(n347) );
  XNOR2_X1 U215 ( .A(n350), .B(n349), .ZN(n294) );
  OR2_X1 U216 ( .A1(n721), .A2(n429), .ZN(n158) );
  NAND2_X1 U217 ( .A1(n183), .A2(n182), .ZN(n471) );
  BUF_X2 U218 ( .A(a_in[9]), .Z(n748) );
  NAND2_X1 U219 ( .A1(n190), .A2(n188), .ZN(n178) );
  OR2_X1 U220 ( .A1(n278), .A2(n195), .ZN(n169) );
  OR2_X1 U221 ( .A1(n447), .A2(n751), .ZN(n445) );
  XNOR2_X1 U222 ( .A(n447), .B(n751), .ZN(n151) );
  NAND2_X1 U223 ( .A1(n447), .A2(n751), .ZN(n448) );
  OR2_X1 U224 ( .A1(n420), .A2(n126), .ZN(n421) );
  NAND2_X1 U225 ( .A1(n542), .A2(n538), .ZN(n539) );
  XOR2_X1 U226 ( .A(n760), .B(a_in[2]), .Z(n174) );
  INV_X1 U227 ( .A(n499), .ZN(n131) );
  NOR2_X1 U228 ( .A1(n498), .A2(n497), .ZN(n546) );
  BUF_X1 U229 ( .A(n291), .Z(n132) );
  BUF_X1 U230 ( .A(n291), .Z(n133) );
  BUF_X1 U231 ( .A(n291), .Z(n423) );
  NOR2_X2 U232 ( .A1(n592), .A2(reset), .ZN(n134) );
  NOR2_X1 U233 ( .A1(n568), .A2(n530), .ZN(n135) );
  OR2_X1 U234 ( .A1(n90), .A2(n116), .ZN(n137) );
  OR2_X1 U235 ( .A1(n393), .A2(n392), .ZN(n143) );
  AND2_X1 U236 ( .A1(n745), .A2(f[18]), .ZN(n144) );
  OR2_X1 U237 ( .A1(n670), .A2(n683), .ZN(n145) );
  AND2_X1 U238 ( .A1(n355), .A2(f[7]), .ZN(n381) );
  AND2_X1 U239 ( .A1(n536), .A2(n789), .ZN(n146) );
  OR2_X1 U240 ( .A1(n560), .A2(n530), .ZN(n147) );
  XNOR2_X1 U244 ( .A(a_in[1]), .B(n771), .ZN(n309) );
  XNOR2_X1 U245 ( .A(n749), .B(b_in[9]), .ZN(n171) );
  OAI22_X1 U246 ( .A1(n344), .A2(n171), .B1(n342), .B2(n104), .ZN(n181) );
  NOR2_X1 U247 ( .A1(n764), .A2(n139), .ZN(n164) );
  XOR2_X1 U248 ( .A(a_in[6]), .B(a_in[7]), .Z(n148) );
  XNOR2_X1 U249 ( .A(n750), .B(a_in[6]), .ZN(n149) );
  NAND2_X1 U250 ( .A1(n148), .A2(n149), .ZN(n194) );
  BUF_X1 U251 ( .A(n194), .Z(n278) );
  BUF_X2 U252 ( .A(a_in[7]), .Z(n417) );
  XNOR2_X1 U253 ( .A(n417), .B(b_in[5]), .ZN(n165) );
  XNOR2_X1 U254 ( .A(n417), .B(b_in[6]), .ZN(n150) );
  OAI22_X1 U255 ( .A1(n278), .A2(n165), .B1(n524), .B2(n150), .ZN(n179) );
  BUF_X1 U256 ( .A(n194), .Z(n484) );
  XNOR2_X1 U257 ( .A(n417), .B(b_in[7]), .ZN(n431) );
  OAI22_X1 U258 ( .A1(n484), .A2(n150), .B1(n524), .B2(n431), .ZN(n447) );
  XNOR2_X1 U259 ( .A(n446), .B(n151), .ZN(n473) );
  XOR2_X1 U260 ( .A(n759), .B(n772), .Z(n152) );
  XNOR2_X1 U261 ( .A(\DP_OP_12J1_122_830/n469 ), .B(a_in[4]), .ZN(n201) );
  NAND2_X1 U262 ( .A1(n152), .A2(n201), .ZN(n291) );
  XNOR2_X1 U263 ( .A(n115), .B(b_in[8]), .ZN(n156) );
  XNOR2_X1 U264 ( .A(n115), .B(b_in[9]), .ZN(n422) );
  BUF_X2 U265 ( .A(n201), .Z(n420) );
  OR2_X1 U266 ( .A1(n422), .A2(n420), .ZN(n153) );
  OAI21_X1 U267 ( .B1(n423), .B2(n156), .A(n153), .ZN(n433) );
  NOR2_X1 U268 ( .A1(n764), .A2(n770), .ZN(n434) );
  XNOR2_X1 U269 ( .A(n433), .B(n154), .ZN(n458) );
  XNOR2_X1 U270 ( .A(n758), .B(n757), .ZN(n205) );
  XNOR2_X1 U271 ( .A(n757), .B(a_in[9]), .ZN(n155) );
  NAND2_X1 U272 ( .A1(n86), .A2(n155), .ZN(n204) );
  BUF_X2 U273 ( .A(a_in[9]), .Z(n487) );
  XNOR2_X1 U274 ( .A(n487), .B(b_in[3]), .ZN(n166) );
  BUF_X2 U275 ( .A(n86), .Z(n721) );
  XNOR2_X1 U276 ( .A(n487), .B(b_in[4]), .ZN(n159) );
  OAI22_X1 U277 ( .A1(n103), .A2(n166), .B1(n721), .B2(n159), .ZN(n211) );
  XNOR2_X1 U278 ( .A(n114), .B(b_in[7]), .ZN(n163) );
  OAI22_X1 U279 ( .A1(n423), .A2(n163), .B1(n420), .B2(n156), .ZN(n210) );
  AND2_X1 U280 ( .A1(a_in[9]), .A2(b_in[2]), .ZN(n157) );
  XNOR2_X1 U281 ( .A(n456), .B(n458), .ZN(n162) );
  AOI21_X1 U282 ( .B1(n344), .B2(n342), .A(n104), .ZN(n443) );
  FA_X1 U283 ( .A(f[12]), .B(n92), .CI(n157), .CO(n440), .S(n209) );
  XNOR2_X1 U284 ( .A(n443), .B(n440), .ZN(n161) );
  XNOR2_X1 U285 ( .A(n487), .B(b_in[5]), .ZN(n429) );
  INV_X1 U286 ( .A(n441), .ZN(n160) );
  XNOR2_X1 U287 ( .A(n161), .B(n160), .ZN(n457) );
  XNOR2_X1 U288 ( .A(n162), .B(n457), .ZN(n472) );
  AND2_X1 U289 ( .A1(b_in[0]), .A2(n487), .ZN(n221) );
  XNOR2_X1 U290 ( .A(n92), .B(b_in[9]), .ZN(n200) );
  OR2_X2 U291 ( .A1(a_in[0]), .A2(n762), .ZN(n358) );
  OAI22_X1 U292 ( .A1(n200), .A2(n358), .B1(n751), .B2(n769), .ZN(n220) );
  XNOR2_X1 U293 ( .A(n114), .B(b_in[6]), .ZN(n196) );
  FA_X1 U294 ( .A(f[11]), .B(n102), .CI(n164), .CO(n180), .S(n227) );
  XNOR2_X1 U295 ( .A(n417), .B(b_in[4]), .ZN(n195) );
  OR2_X1 U296 ( .A1(n165), .A2(n524), .ZN(n168) );
  NAND2_X1 U297 ( .A1(n169), .A2(n168), .ZN(n190) );
  XNOR2_X1 U298 ( .A(n487), .B(b_in[2]), .ZN(n192) );
  OAI22_X1 U299 ( .A1(n103), .A2(n192), .B1(n721), .B2(n166), .ZN(n188) );
  INV_X1 U300 ( .A(n188), .ZN(n167) );
  AND2_X1 U301 ( .A1(n168), .A2(n167), .ZN(n170) );
  NAND2_X1 U302 ( .A1(n170), .A2(n169), .ZN(n176) );
  XNOR2_X1 U303 ( .A(n749), .B(b_in[8]), .ZN(n193) );
  OR2_X1 U304 ( .A1(n117), .A2(n193), .ZN(n175) );
  INV_X1 U305 ( .A(n171), .ZN(n172) );
  NAND2_X1 U306 ( .A1(n172), .A2(n117), .ZN(n173) );
  OAI21_X1 U307 ( .B1(n175), .B2(n174), .A(n173), .ZN(n189) );
  NAND2_X1 U308 ( .A1(n176), .A2(n124), .ZN(n177) );
  NAND2_X1 U309 ( .A1(n178), .A2(n177), .ZN(n184) );
  FA_X1 U310 ( .A(n181), .B(n180), .CI(n179), .CO(n446), .S(n186) );
  OAI21_X1 U311 ( .B1(n185), .B2(n184), .A(n186), .ZN(n183) );
  NAND2_X1 U312 ( .A1(n185), .A2(n184), .ZN(n182) );
  XNOR2_X1 U313 ( .A(n185), .B(n85), .ZN(n187) );
  XNOR2_X1 U314 ( .A(n187), .B(n186), .ZN(n255) );
  XNOR2_X1 U315 ( .A(n188), .B(n189), .ZN(n191) );
  XNOR2_X1 U316 ( .A(n191), .B(n190), .ZN(n232) );
  XNOR2_X1 U317 ( .A(n748), .B(b_in[1]), .ZN(n197) );
  OAI22_X1 U318 ( .A1(n722), .A2(n197), .B1(n721), .B2(n192), .ZN(n219) );
  XNOR2_X1 U319 ( .A(n96), .B(b_in[7]), .ZN(n223) );
  OAI22_X1 U320 ( .A1(n113), .A2(n223), .B1(n342), .B2(n193), .ZN(n218) );
  BUF_X1 U321 ( .A(n194), .Z(n418) );
  XNOR2_X1 U322 ( .A(n417), .B(b_in[3]), .ZN(n222) );
  OAI22_X1 U323 ( .A1(n418), .A2(n222), .B1(n524), .B2(n195), .ZN(n217) );
  XNOR2_X1 U324 ( .A(n114), .B(b_in[5]), .ZN(n202) );
  OAI22_X1 U325 ( .A1(n133), .A2(n202), .B1(n420), .B2(n196), .ZN(n242) );
  XNOR2_X1 U326 ( .A(n748), .B(b_in[0]), .ZN(n199) );
  OR2_X1 U327 ( .A1(n205), .A2(n197), .ZN(n198) );
  OAI21_X1 U328 ( .B1(n722), .B2(n199), .A(n198), .ZN(n224) );
  XNOR2_X1 U329 ( .A(n335), .B(n91), .ZN(n238) );
  OAI22_X1 U330 ( .A1(n238), .A2(n358), .B1(n200), .B2(n769), .ZN(n241) );
  XNOR2_X1 U331 ( .A(n115), .B(b_in[4]), .ZN(n235) );
  INV_X1 U332 ( .A(n201), .ZN(n292) );
  INV_X1 U333 ( .A(n292), .ZN(n203) );
  OAI22_X1 U334 ( .A1(n235), .A2(n291), .B1(n203), .B2(n202), .ZN(n240) );
  OR2_X1 U335 ( .A1(b_in[0]), .A2(n764), .ZN(n206) );
  OAI22_X1 U336 ( .A1(n103), .A2(n764), .B1(n721), .B2(n206), .ZN(n239) );
  OAI21_X1 U337 ( .B1(n242), .B2(n243), .A(n244), .ZN(n208) );
  NAND2_X1 U338 ( .A1(n243), .A2(n242), .ZN(n207) );
  NAND2_X1 U339 ( .A1(n208), .A2(n207), .ZN(n230) );
  INV_X1 U340 ( .A(n254), .ZN(n213) );
  FA_X1 U341 ( .A(n209), .B(n211), .CI(n210), .CO(n456), .S(n253) );
  INV_X1 U342 ( .A(n253), .ZN(n212) );
  NAND2_X1 U343 ( .A1(n213), .A2(n212), .ZN(n214) );
  NAND2_X1 U344 ( .A1(n214), .A2(n255), .ZN(n216) );
  NAND2_X1 U345 ( .A1(n106), .A2(n253), .ZN(n215) );
  NAND2_X1 U346 ( .A1(n216), .A2(n215), .ZN(n414) );
  NOR2_X1 U347 ( .A1(n415), .A2(n123), .ZN(n416) );
  FA_X1 U348 ( .A(n219), .B(n218), .CI(n217), .CO(n231), .S(n246) );
  FA_X1 U349 ( .A(n221), .B(f[10]), .CI(n220), .CO(n229), .S(n247) );
  XNOR2_X1 U350 ( .A(n417), .B(n111), .ZN(n234) );
  OAI22_X1 U351 ( .A1(n418), .A2(n234), .B1(n524), .B2(n222), .ZN(n284) );
  XNOR2_X1 U352 ( .A(n96), .B(b_in[6]), .ZN(n237) );
  OAI22_X1 U353 ( .A1(n113), .A2(n237), .B1(n342), .B2(n223), .ZN(n283) );
  XNOR2_X1 U354 ( .A(n224), .B(n763), .ZN(n282) );
  OAI21_X1 U355 ( .B1(n246), .B2(n247), .A(n248), .ZN(n226) );
  NAND2_X1 U356 ( .A1(n246), .A2(n247), .ZN(n225) );
  NAND2_X1 U357 ( .A1(n226), .A2(n225), .ZN(n257) );
  XNOR2_X1 U358 ( .A(n257), .B(n262), .ZN(n233) );
  FA_X1 U359 ( .A(n232), .B(n231), .CI(n230), .CO(n254), .S(n260) );
  XNOR2_X1 U360 ( .A(n233), .B(n260), .ZN(n577) );
  XNOR2_X1 U361 ( .A(n417), .B(b_in[1]), .ZN(n276) );
  OAI22_X1 U362 ( .A1(n484), .A2(n276), .B1(n524), .B2(n234), .ZN(n379) );
  XNOR2_X1 U363 ( .A(n114), .B(b_in[3]), .ZN(n272) );
  OR2_X1 U364 ( .A1(n420), .A2(n235), .ZN(n236) );
  OAI21_X1 U365 ( .B1(n133), .B2(n272), .A(n236), .ZN(n378) );
  XNOR2_X1 U366 ( .A(n96), .B(b_in[5]), .ZN(n273) );
  OAI22_X1 U367 ( .A1(n113), .A2(n273), .B1(n342), .B2(n237), .ZN(n377) );
  OAI22_X1 U368 ( .A1(n358), .A2(n356), .B1(n238), .B2(n769), .ZN(n274) );
  FA_X1 U369 ( .A(n241), .B(n240), .CI(n239), .CO(n244), .S(n268) );
  XNOR2_X1 U370 ( .A(n248), .B(n247), .ZN(n249) );
  XNOR2_X1 U371 ( .A(n249), .B(n250), .ZN(n266) );
  OAI21_X1 U372 ( .B1(n265), .B2(n264), .A(n266), .ZN(n252) );
  NAND2_X1 U373 ( .A1(n265), .A2(n264), .ZN(n251) );
  NAND2_X1 U374 ( .A1(n252), .A2(n251), .ZN(n576) );
  NOR2_X1 U375 ( .A1(n577), .A2(n576), .ZN(n409) );
  NOR2_X1 U376 ( .A1(n416), .A2(n409), .ZN(n288) );
  XNOR2_X1 U377 ( .A(n254), .B(n253), .ZN(n256) );
  XNOR2_X1 U378 ( .A(n256), .B(n255), .ZN(n578) );
  INV_X1 U379 ( .A(n257), .ZN(n261) );
  NAND2_X1 U380 ( .A1(n261), .A2(n258), .ZN(n259) );
  NAND2_X1 U381 ( .A1(n259), .A2(n260), .ZN(n412) );
  INV_X1 U382 ( .A(n261), .ZN(n263) );
  NAND2_X1 U383 ( .A1(n263), .A2(n262), .ZN(n411) );
  NOR2_X1 U384 ( .A1(n578), .A2(n413), .ZN(n410) );
  XNOR2_X1 U385 ( .A(n265), .B(n264), .ZN(n267) );
  XNOR2_X1 U386 ( .A(n267), .B(n266), .ZN(n408) );
  FA_X1 U387 ( .A(n268), .B(n269), .CI(n270), .CO(n265), .S(n399) );
  INV_X1 U388 ( .A(n417), .ZN(n523) );
  OR2_X1 U389 ( .A1(b_in[0]), .A2(n523), .ZN(n271) );
  OAI22_X1 U390 ( .A1(n418), .A2(n523), .B1(n271), .B2(n524), .ZN(n363) );
  XNOR2_X1 U391 ( .A(n115), .B(n111), .ZN(n345) );
  OAI22_X1 U392 ( .A1(n132), .A2(n345), .B1(n420), .B2(n272), .ZN(n362) );
  XNOR2_X1 U393 ( .A(n749), .B(b_in[4]), .ZN(n341) );
  OAI22_X1 U394 ( .A1(n113), .A2(n341), .B1(n342), .B2(n273), .ZN(n361) );
  FA_X1 U395 ( .A(n275), .B(f[8]), .CI(n274), .CO(n269), .S(n380) );
  XNOR2_X1 U396 ( .A(n417), .B(n108), .ZN(n277) );
  OAI22_X1 U397 ( .A1(n278), .A2(n277), .B1(n524), .B2(n276), .ZN(n355) );
  OR2_X1 U398 ( .A1(n381), .A2(n380), .ZN(n279) );
  NAND2_X1 U399 ( .A1(n382), .A2(n279), .ZN(n281) );
  NAND2_X1 U400 ( .A1(n381), .A2(n125), .ZN(n280) );
  FA_X1 U401 ( .A(n284), .B(n283), .CI(n282), .CO(n248), .S(n392) );
  NAND2_X1 U402 ( .A1(n393), .A2(n392), .ZN(n285) );
  NOR2_X1 U403 ( .A1(n410), .A2(n670), .ZN(n287) );
  XNOR2_X1 U404 ( .A(n749), .B(n111), .ZN(n297) );
  XNOR2_X1 U405 ( .A(n749), .B(b_in[3]), .ZN(n343) );
  OAI22_X1 U406 ( .A1(n113), .A2(n297), .B1(n342), .B2(n343), .ZN(n339) );
  XNOR2_X1 U407 ( .A(n92), .B(b_in[4]), .ZN(n293) );
  OAI22_X1 U408 ( .A1(n358), .A2(n293), .B1(n336), .B2(n769), .ZN(n338) );
  OR2_X1 U409 ( .A1(b_in[0]), .A2(n126), .ZN(n289) );
  OAI22_X1 U410 ( .A1(n132), .A2(n126), .B1(n289), .B2(n420), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n114), .B(b_in[0]), .ZN(n290) );
  XNOR2_X1 U412 ( .A(n115), .B(b_in[1]), .ZN(n346) );
  OAI22_X1 U413 ( .A1(n290), .A2(n291), .B1(n203), .B2(n346), .ZN(n340) );
  AND2_X1 U414 ( .A1(n292), .A2(b_in[0]), .ZN(n296) );
  XNOR2_X1 U415 ( .A(n762), .B(n770), .ZN(n298) );
  OAI22_X1 U416 ( .A1(n358), .A2(n298), .B1(n293), .B2(n769), .ZN(n295) );
  FA_X1 U417 ( .A(n296), .B(f[4]), .CI(n295), .CO(n349), .S(n325) );
  XNOR2_X1 U418 ( .A(n749), .B(b_in[1]), .ZN(n306) );
  OAI22_X1 U419 ( .A1(n344), .A2(n306), .B1(n342), .B2(n297), .ZN(n324) );
  INV_X1 U420 ( .A(n324), .ZN(n301) );
  XNOR2_X1 U421 ( .A(n92), .B(b_in[2]), .ZN(n299) );
  OAI22_X1 U422 ( .A1(n358), .A2(n299), .B1(n298), .B2(n769), .ZN(n308) );
  INV_X1 U423 ( .A(n323), .ZN(n300) );
  NAND2_X1 U424 ( .A1(n301), .A2(n300), .ZN(n302) );
  NAND2_X1 U425 ( .A1(n325), .A2(n302), .ZN(n304) );
  NAND2_X1 U426 ( .A1(n324), .A2(n323), .ZN(n303) );
  NAND2_X1 U427 ( .A1(n304), .A2(n303), .ZN(n333) );
  NOR2_X1 U428 ( .A1(n334), .A2(n333), .ZN(n636) );
  OR2_X1 U429 ( .A1(b_in[0]), .A2(n104), .ZN(n305) );
  OAI22_X1 U430 ( .A1(n113), .A2(n104), .B1(n305), .B2(n342), .ZN(n329) );
  XNOR2_X1 U431 ( .A(n96), .B(b_in[0]), .ZN(n307) );
  OAI22_X1 U432 ( .A1(n113), .A2(n307), .B1(n342), .B2(n306), .ZN(n328) );
  HA_X1 U433 ( .A(n308), .B(f[3]), .CO(n323), .S(n327) );
  AND2_X1 U434 ( .A1(b_in[0]), .A2(n117), .ZN(n312) );
  XNOR2_X1 U435 ( .A(n335), .B(b_in[1]), .ZN(n313) );
  XNOR2_X1 U436 ( .A(n92), .B(b_in[2]), .ZN(n310) );
  OAI22_X1 U437 ( .A1(n313), .A2(n358), .B1(n310), .B2(n769), .ZN(n311) );
  NOR2_X1 U438 ( .A1(n321), .A2(n320), .ZN(n620) );
  FA_X1 U439 ( .A(n312), .B(f[2]), .CI(n311), .CO(n320), .S(n319) );
  OAI22_X1 U440 ( .A1(n358), .A2(b_in[0]), .B1(n313), .B2(n769), .ZN(n314) );
  OR2_X1 U441 ( .A1(n318), .A2(n319), .ZN(n624) );
  HA_X1 U442 ( .A(n314), .B(f[1]), .CO(n318), .S(n317) );
  OR2_X1 U443 ( .A1(n108), .A2(n751), .ZN(n315) );
  NAND2_X1 U444 ( .A1(n315), .A2(n358), .ZN(n316) );
  NOR2_X1 U445 ( .A1(n317), .A2(n316), .ZN(n603) );
  AND2_X1 U446 ( .A1(n108), .A2(a_in[0]), .ZN(n593) );
  NAND2_X1 U447 ( .A1(n593), .A2(f[0]), .ZN(n606) );
  NAND2_X1 U448 ( .A1(n317), .A2(n316), .ZN(n604) );
  AOI21_X1 U449 ( .B1(n624), .B2(n623), .A(n95), .ZN(n322) );
  NAND2_X1 U450 ( .A1(n321), .A2(n320), .ZN(n621) );
  OAI21_X1 U451 ( .B1(n620), .B2(n322), .A(n621), .ZN(n616) );
  FA_X1 U452 ( .A(n329), .B(n328), .CI(n327), .CO(n330), .S(n321) );
  OR2_X1 U453 ( .A1(n331), .A2(n330), .ZN(n615) );
  NAND2_X1 U454 ( .A1(n331), .A2(n330), .ZN(n614) );
  INV_X1 U455 ( .A(n614), .ZN(n332) );
  AOI21_X1 U456 ( .B1(n616), .B2(n615), .A(n332), .ZN(n635) );
  NAND2_X1 U457 ( .A1(n334), .A2(n333), .ZN(n637) );
  OAI21_X1 U458 ( .B1(n635), .B2(n636), .A(n637), .ZN(n645) );
  XNOR2_X1 U459 ( .A(n102), .B(b_in[6]), .ZN(n357) );
  OAI22_X1 U460 ( .A1(n336), .A2(n358), .B1(n357), .B2(n769), .ZN(n360) );
  NOR2_X1 U461 ( .A1(n761), .A2(n524), .ZN(n359) );
  FA_X1 U462 ( .A(n339), .B(n338), .CI(n337), .CO(n369), .S(n348) );
  HA_X1 U463 ( .A(n340), .B(f[5]), .CO(n366), .S(n350) );
  OAI22_X1 U464 ( .A1(n344), .A2(n343), .B1(n342), .B2(n341), .ZN(n365) );
  OAI22_X1 U465 ( .A1(n132), .A2(n346), .B1(n420), .B2(n345), .ZN(n364) );
  AOI21_X1 U466 ( .B1(n645), .B2(n644), .A(n643), .ZN(n373) );
  XNOR2_X1 U467 ( .A(n355), .B(n756), .ZN(n376) );
  OAI22_X1 U468 ( .A1(n358), .A2(n357), .B1(n356), .B2(n769), .ZN(n375) );
  FA_X1 U469 ( .A(n360), .B(f[6]), .CI(n359), .CO(n374), .S(n370) );
  FA_X1 U470 ( .A(n363), .B(n362), .CI(n361), .CO(n382), .S(n389) );
  FA_X1 U471 ( .A(n364), .B(n365), .CI(n366), .CO(n388), .S(n368) );
  XNOR2_X1 U472 ( .A(n389), .B(n388), .ZN(n367) );
  FA_X1 U473 ( .A(n370), .B(n369), .CI(n368), .CO(n371), .S(n354) );
  NOR2_X1 U474 ( .A1(n372), .A2(n371), .ZN(n647) );
  NAND2_X1 U475 ( .A1(n372), .A2(n371), .ZN(n648) );
  OAI21_X1 U476 ( .B1(n373), .B2(n647), .A(n648), .ZN(n653) );
  FA_X1 U477 ( .A(n376), .B(n375), .CI(n374), .CO(n396), .S(n386) );
  FA_X1 U478 ( .A(n379), .B(n378), .CI(n377), .CO(n270), .S(n395) );
  XNOR2_X1 U479 ( .A(n380), .B(n381), .ZN(n383) );
  XNOR2_X1 U480 ( .A(n383), .B(n382), .ZN(n394) );
  NAND2_X1 U481 ( .A1(n387), .A2(n386), .ZN(n391) );
  NAND2_X1 U482 ( .A1(n391), .A2(n390), .ZN(n402) );
  NOR2_X1 U483 ( .A1(n403), .A2(n402), .ZN(n655) );
  XNOR2_X1 U484 ( .A(n93), .B(n392), .ZN(n400) );
  XNOR2_X1 U485 ( .A(n399), .B(n400), .ZN(n405) );
  FA_X1 U486 ( .A(n396), .B(n395), .CI(n394), .CO(n404), .S(n403) );
  NOR2_X1 U487 ( .A1(n404), .A2(n405), .ZN(n397) );
  NOR2_X1 U488 ( .A1(n397), .A2(n655), .ZN(n398) );
  NAND2_X1 U489 ( .A1(n653), .A2(n398), .ZN(n575) );
  XNOR2_X1 U490 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U491 ( .A1(n401), .A2(n404), .ZN(n664) );
  NAND2_X1 U492 ( .A1(n403), .A2(n402), .ZN(n657) );
  NAND2_X1 U493 ( .A1(n405), .A2(n404), .ZN(n665) );
  OAI21_X1 U494 ( .B1(n664), .B2(n657), .A(n665), .ZN(n406) );
  INV_X1 U495 ( .A(n406), .ZN(n574) );
  NAND2_X1 U496 ( .A1(n575), .A2(n574), .ZN(n700) );
  NAND2_X1 U497 ( .A1(n700), .A2(n701), .ZN(n513) );
  NAND2_X1 U498 ( .A1(n408), .A2(n407), .ZN(n671) );
  NAND2_X1 U499 ( .A1(n121), .A2(n576), .ZN(n684) );
  OAI21_X1 U500 ( .B1(n409), .B2(n671), .A(n684), .ZN(n580) );
  NOR2_X1 U501 ( .A1(n415), .A2(n123), .ZN(n585) );
  NOR2_X1 U502 ( .A1(n585), .A2(n410), .ZN(n544) );
  NAND2_X1 U503 ( .A1(n412), .A2(n411), .ZN(n413) );
  NAND2_X1 U504 ( .A1(n90), .A2(n116), .ZN(n693) );
  NAND2_X1 U505 ( .A1(n415), .A2(n414), .ZN(n586) );
  OAI21_X1 U506 ( .B1(n110), .B2(n693), .A(n586), .ZN(n543) );
  AOI21_X1 U507 ( .B1(n580), .B2(n544), .A(n543), .ZN(n512) );
  XNOR2_X1 U508 ( .A(n417), .B(b_in[8]), .ZN(n430) );
  XNOR2_X1 U509 ( .A(n417), .B(b_in[9]), .ZN(n485) );
  OAI22_X1 U510 ( .A1(n418), .A2(n430), .B1(n524), .B2(n485), .ZN(n491) );
  XNOR2_X1 U511 ( .A(n748), .B(b_in[6]), .ZN(n428) );
  XNOR2_X1 U512 ( .A(n487), .B(b_in[7]), .ZN(n488) );
  OAI22_X1 U513 ( .A1(n122), .A2(n428), .B1(n721), .B2(n488), .ZN(n490) );
  AOI21_X1 U514 ( .B1(n132), .B2(n420), .A(n126), .ZN(n419) );
  INV_X1 U515 ( .A(n419), .ZN(n489) );
  OAI21_X1 U516 ( .B1(n133), .B2(n422), .A(n421), .ZN(n439) );
  NOR2_X1 U517 ( .A1(n764), .A2(n140), .ZN(n437) );
  NAND2_X1 U518 ( .A1(n439), .A2(n424), .ZN(n426) );
  NAND2_X1 U519 ( .A1(n426), .A2(n425), .ZN(n481) );
  NOR2_X1 U520 ( .A1(n764), .A2(n768), .ZN(n486) );
  XNOR2_X1 U521 ( .A(n481), .B(n480), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n479), .B(n427), .ZN(n492) );
  OAI22_X1 U523 ( .A1(n103), .A2(n429), .B1(n128), .B2(n428), .ZN(n463) );
  OAI22_X1 U524 ( .A1(n484), .A2(n431), .B1(n524), .B2(n430), .ZN(n462) );
  NAND2_X1 U525 ( .A1(n433), .A2(n432), .ZN(n436) );
  XNOR2_X1 U526 ( .A(n492), .B(n493), .ZN(n455) );
  XNOR2_X1 U527 ( .A(n439), .B(n438), .ZN(n465) );
  AND2_X1 U528 ( .A1(n465), .A2(n464), .ZN(n453) );
  NAND2_X1 U529 ( .A1(n446), .A2(n445), .ZN(n449) );
  NAND2_X1 U530 ( .A1(n449), .A2(n448), .ZN(n467) );
  INV_X1 U531 ( .A(n465), .ZN(n451) );
  INV_X1 U532 ( .A(n464), .ZN(n450) );
  NAND2_X1 U533 ( .A1(n451), .A2(n450), .ZN(n452) );
  OAI21_X1 U534 ( .B1(n453), .B2(n467), .A(n452), .ZN(n454) );
  INV_X1 U535 ( .A(n454), .ZN(n494) );
  XNOR2_X1 U536 ( .A(n455), .B(n494), .ZN(n475) );
  OAI21_X1 U537 ( .B1(n457), .B2(n458), .A(n456), .ZN(n460) );
  NAND2_X1 U538 ( .A1(n457), .A2(n458), .ZN(n459) );
  NAND2_X1 U539 ( .A1(n460), .A2(n459), .ZN(n470) );
  FA_X1 U540 ( .A(n463), .B(n462), .CI(n461), .CO(n493), .S(n469) );
  XNOR2_X1 U541 ( .A(n464), .B(n465), .ZN(n466) );
  XNOR2_X1 U542 ( .A(n467), .B(n466), .ZN(n468) );
  FA_X1 U543 ( .A(n470), .B(n469), .CI(n468), .CO(n474), .S(n501) );
  FA_X1 U544 ( .A(n472), .B(n473), .CI(n471), .CO(n676), .S(n415) );
  NAND2_X1 U545 ( .A1(n501), .A2(n676), .ZN(n702) );
  NAND2_X1 U546 ( .A1(n475), .A2(n474), .ZN(n707) );
  OAI21_X1 U547 ( .B1(n706), .B2(n702), .A(n707), .ZN(n566) );
  NAND3_X1 U548 ( .A1(n129), .A2(n512), .A3(n532), .ZN(n511) );
  INV_X1 U549 ( .A(n481), .ZN(n477) );
  NAND2_X1 U550 ( .A1(n479), .A2(n478), .ZN(n483) );
  NOR2_X1 U551 ( .A1(n764), .A2(n767), .ZN(n522) );
  OAI22_X1 U552 ( .A1(n525), .A2(n485), .B1(n524), .B2(n523), .ZN(n521) );
  FA_X1 U553 ( .A(f[15]), .B(f[14]), .CI(n486), .CO(n520), .S(n480) );
  XNOR2_X1 U554 ( .A(n487), .B(b_in[8]), .ZN(n527) );
  OAI22_X1 U555 ( .A1(n103), .A2(n488), .B1(n128), .B2(n527), .ZN(n519) );
  FA_X1 U556 ( .A(n491), .B(n490), .CI(n489), .CO(n518), .S(n479) );
  INV_X1 U557 ( .A(n546), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n498), .A2(n497), .ZN(n563) );
  AND2_X1 U559 ( .A1(n499), .A2(n563), .ZN(n500) );
  INV_X1 U560 ( .A(n500), .ZN(n503) );
  NOR2_X2 U561 ( .A1(n773), .A2(reset), .ZN(n789) );
  INV_X1 U562 ( .A(n789), .ZN(n530) );
  OR2_X1 U563 ( .A1(n503), .A2(n530), .ZN(n510) );
  BUF_X1 U564 ( .A(n501), .Z(n677) );
  NOR2_X1 U565 ( .A1(n677), .A2(n676), .ZN(n502) );
  NOR2_X1 U566 ( .A1(n502), .A2(n706), .ZN(n547) );
  NAND2_X1 U567 ( .A1(n532), .A2(n89), .ZN(n506) );
  NOR2_X2 U568 ( .A1(enable_f), .A2(reset), .ZN(n745) );
  NAND2_X1 U569 ( .A1(n745), .A2(f[16]), .ZN(n505) );
  OAI21_X1 U570 ( .B1(n510), .B2(n506), .A(n505), .ZN(n507) );
  INV_X1 U571 ( .A(n507), .ZN(n508) );
  OAI211_X1 U572 ( .C1(n511), .C2(n510), .A(n509), .B(n508), .ZN(n48) );
  NAND2_X1 U573 ( .A1(n513), .A2(n512), .ZN(n679) );
  NOR2_X1 U574 ( .A1(n89), .A2(n131), .ZN(n514) );
  NAND2_X1 U575 ( .A1(n679), .A2(n514), .ZN(n542) );
  FA_X1 U576 ( .A(n517), .B(n516), .CI(n515), .CO(n529), .S(n498) );
  FA_X1 U577 ( .A(n520), .B(n519), .CI(n518), .CO(n551), .S(n515) );
  FA_X1 U578 ( .A(n522), .B(n138), .CI(n521), .CO(n550), .S(n516) );
  AOI21_X1 U579 ( .B1(n525), .B2(n524), .A(n523), .ZN(n526) );
  INV_X1 U580 ( .A(n526), .ZN(n556) );
  XNOR2_X1 U581 ( .A(n748), .B(b_in[9]), .ZN(n552) );
  OAI22_X1 U582 ( .A1(n722), .A2(n527), .B1(n128), .B2(n552), .ZN(n555) );
  NOR2_X1 U583 ( .A1(n764), .A2(n766), .ZN(n553) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n561) );
  AND2_X1 U585 ( .A1(n120), .A2(n561), .ZN(n536) );
  INV_X1 U586 ( .A(n105), .ZN(n532) );
  OAI21_X1 U587 ( .B1(n532), .B2(n131), .A(n563), .ZN(n533) );
  INV_X1 U588 ( .A(n533), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n745), .A2(f[17]), .ZN(n534) );
  OAI211_X1 U590 ( .C1(n542), .C2(n541), .A(n540), .B(n539), .ZN(n47) );
  AOI21_X1 U591 ( .B1(n580), .B2(n544), .A(n543), .ZN(n705) );
  NAND2_X1 U592 ( .A1(n700), .A2(n701), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n545), .A2(n705), .ZN(n734) );
  NOR2_X1 U594 ( .A1(n546), .A2(n119), .ZN(n565) );
  NAND2_X1 U595 ( .A1(n565), .A2(n547), .ZN(n732) );
  INV_X1 U596 ( .A(n732), .ZN(n548) );
  AND2_X1 U597 ( .A1(n734), .A2(n548), .ZN(n569) );
  FA_X1 U598 ( .A(n551), .B(n550), .CI(n549), .CO(n558), .S(n528) );
  NOR2_X1 U599 ( .A1(n764), .A2(n141), .ZN(n720) );
  OAI22_X1 U600 ( .A1(n122), .A2(n552), .B1(n128), .B2(n764), .ZN(n719) );
  FA_X1 U601 ( .A(f[17]), .B(f[16]), .CI(n553), .CO(n715), .S(n554) );
  FA_X1 U602 ( .A(n556), .B(n555), .CI(n554), .CO(n714), .S(n549) );
  NOR2_X1 U603 ( .A1(n558), .A2(n557), .ZN(n736) );
  INV_X1 U604 ( .A(n736), .ZN(n559) );
  NAND2_X1 U605 ( .A1(n558), .A2(n557), .ZN(n735) );
  AND2_X1 U606 ( .A1(n559), .A2(n735), .ZN(n568) );
  OR2_X1 U607 ( .A1(n569), .A2(n147), .ZN(n573) );
  OAI21_X1 U608 ( .B1(n563), .B2(n562), .A(n561), .ZN(n564) );
  AOI21_X1 U609 ( .B1(n565), .B2(n566), .A(n564), .ZN(n737) );
  INV_X1 U610 ( .A(n567), .ZN(n572) );
  AOI21_X1 U611 ( .B1(n569), .B2(n135), .A(n144), .ZN(n571) );
  NAND2_X1 U612 ( .A1(n572), .A2(n135), .ZN(n570) );
  OAI211_X1 U613 ( .C1(n573), .C2(n572), .A(n571), .B(n570), .ZN(n46) );
  AND2_X1 U614 ( .A1(n575), .A2(n574), .ZN(n692) );
  INV_X1 U615 ( .A(n692), .ZN(n674) );
  NOR2_X1 U616 ( .A1(n121), .A2(n576), .ZN(n683) );
  INV_X1 U617 ( .A(n137), .ZN(n581) );
  NOR2_X1 U618 ( .A1(n145), .A2(n581), .ZN(n579) );
  NAND2_X1 U619 ( .A1(n674), .A2(n579), .ZN(n584) );
  INV_X1 U620 ( .A(n580), .ZN(n691) );
  OAI21_X1 U621 ( .B1(n691), .B2(n581), .A(n118), .ZN(n582) );
  INV_X1 U622 ( .A(n582), .ZN(n583) );
  NAND2_X1 U623 ( .A1(n584), .A2(n583), .ZN(n589) );
  INV_X1 U624 ( .A(n585), .ZN(n587) );
  AND2_X1 U625 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U626 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U627 ( .A1(n745), .A2(f[13]), .ZN(n590) );
  OAI21_X1 U628 ( .B1(n591), .B2(n530), .A(n590), .ZN(n51) );
  INV_X1 U629 ( .A(valid_in), .ZN(n592) );
  OR2_X1 U630 ( .A1(n593), .A2(f[0]), .ZN(n594) );
  AND2_X1 U631 ( .A1(n594), .A2(n606), .ZN(n595) );
  AOI22_X1 U632 ( .A1(n595), .A2(n789), .B1(n745), .B2(f[0]), .ZN(n596) );
  INV_X1 U633 ( .A(n596), .ZN(n64) );
  NOR2_X2 U634 ( .A1(valid_in), .A2(reset), .ZN(n752) );
  AOI22_X1 U635 ( .A1(n134), .A2(b[2]), .B1(n752), .B2(n111), .ZN(n787) );
  AOI22_X1 U636 ( .A1(n134), .A2(a[2]), .B1(n752), .B2(a_in[2]), .ZN(n782) );
  AOI22_X1 U637 ( .A1(n134), .A2(b[5]), .B1(n752), .B2(b_in[5]), .ZN(n785) );
  AOI22_X1 U638 ( .A1(n134), .A2(a[8]), .B1(n752), .B2(a_in[8]), .ZN(n779) );
  AOI22_X1 U639 ( .A1(n134), .A2(b[3]), .B1(n752), .B2(b_in[3]), .ZN(n786) );
  AOI22_X1 U640 ( .A1(n134), .A2(b[1]), .B1(n752), .B2(b_in[1]), .ZN(n597) );
  INV_X1 U641 ( .A(n597), .ZN(n73) );
  AOI22_X1 U642 ( .A1(n134), .A2(b[0]), .B1(n752), .B2(n108), .ZN(n598) );
  INV_X1 U643 ( .A(n598), .ZN(n84) );
  AOI22_X1 U644 ( .A1(n134), .A2(b[7]), .B1(n752), .B2(b_in[7]), .ZN(n784) );
  AOI22_X1 U645 ( .A1(n134), .A2(b[4]), .B1(n752), .B2(b_in[4]), .ZN(n599) );
  INV_X1 U646 ( .A(n599), .ZN(n70) );
  AOI22_X1 U647 ( .A1(n134), .A2(b[6]), .B1(n752), .B2(b_in[6]), .ZN(n600) );
  INV_X1 U648 ( .A(n600), .ZN(n68) );
  AOI22_X1 U649 ( .A1(n134), .A2(a[0]), .B1(n752), .B2(a_in[0]), .ZN(n783) );
  AOI22_X1 U650 ( .A1(n134), .A2(a[4]), .B1(n752), .B2(n112), .ZN(n781) );
  AOI22_X1 U651 ( .A1(n134), .A2(a[6]), .B1(n752), .B2(a_in[6]), .ZN(n780) );
  AOI22_X1 U652 ( .A1(n134), .A2(b[8]), .B1(n752), .B2(b_in[8]), .ZN(n601) );
  INV_X1 U653 ( .A(n601), .ZN(n66) );
  AOI22_X1 U654 ( .A1(n134), .A2(b[9]), .B1(n752), .B2(b_in[9]), .ZN(n602) );
  INV_X1 U655 ( .A(n602), .ZN(n65) );
  INV_X1 U656 ( .A(n603), .ZN(n605) );
  NAND2_X1 U657 ( .A1(n605), .A2(n604), .ZN(n607) );
  XOR2_X1 U658 ( .A(n607), .B(n606), .Z(n608) );
  AOI22_X1 U659 ( .A1(n608), .A2(n789), .B1(n745), .B2(f[1]), .ZN(n609) );
  INV_X1 U660 ( .A(n609), .ZN(n63) );
  NAND2_X1 U661 ( .A1(n624), .A2(n610), .ZN(n611) );
  XNOR2_X1 U662 ( .A(n611), .B(n623), .ZN(n612) );
  AOI22_X1 U663 ( .A1(n612), .A2(n789), .B1(n745), .B2(f[2]), .ZN(n613) );
  INV_X1 U664 ( .A(n613), .ZN(n62) );
  NAND2_X1 U665 ( .A1(n615), .A2(n614), .ZN(n617) );
  XNOR2_X1 U666 ( .A(n617), .B(n130), .ZN(n618) );
  AOI22_X1 U667 ( .A1(n618), .A2(n789), .B1(n745), .B2(f[4]), .ZN(n619) );
  INV_X1 U668 ( .A(n619), .ZN(n60) );
  INV_X1 U669 ( .A(n97), .ZN(n622) );
  NAND2_X1 U670 ( .A1(n622), .A2(n621), .ZN(n626) );
  AOI21_X1 U671 ( .B1(n624), .B2(n623), .A(n95), .ZN(n625) );
  XOR2_X1 U672 ( .A(n626), .B(n625), .Z(n627) );
  AOI22_X1 U673 ( .A1(n627), .A2(n789), .B1(n745), .B2(f[3]), .ZN(n628) );
  INV_X1 U674 ( .A(n628), .ZN(n61) );
  NAND2_X1 U675 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U676 ( .A(n632), .B(n631), .ZN(n633) );
  AOI22_X1 U677 ( .A1(n633), .A2(n789), .B1(n745), .B2(f[6]), .ZN(n634) );
  INV_X1 U678 ( .A(n634), .ZN(n58) );
  INV_X1 U679 ( .A(n636), .ZN(n638) );
  NAND2_X1 U680 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U681 ( .A(n640), .B(n639), .Z(n641) );
  AOI22_X1 U682 ( .A1(n641), .A2(n789), .B1(n745), .B2(f[5]), .ZN(n642) );
  INV_X1 U683 ( .A(n642), .ZN(n59) );
  AOI21_X1 U684 ( .B1(n645), .B2(n630), .A(n94), .ZN(n646) );
  INV_X1 U685 ( .A(n647), .ZN(n649) );
  NAND2_X1 U686 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U687 ( .A(n646), .B(n650), .Z(n651) );
  AOI22_X1 U688 ( .A1(n651), .A2(n789), .B1(n745), .B2(f[7]), .ZN(n652) );
  INV_X1 U689 ( .A(n652), .ZN(n57) );
  INV_X1 U690 ( .A(n654), .ZN(n663) );
  INV_X1 U691 ( .A(n656), .ZN(n661) );
  NAND2_X1 U692 ( .A1(n661), .A2(n662), .ZN(n658) );
  XOR2_X1 U693 ( .A(n663), .B(n658), .Z(n659) );
  AOI22_X1 U694 ( .A1(n659), .A2(n789), .B1(n745), .B2(f[8]), .ZN(n660) );
  INV_X1 U695 ( .A(n660), .ZN(n56) );
  OAI21_X1 U696 ( .B1(n663), .B2(n656), .A(n662), .ZN(n667) );
  NAND2_X1 U697 ( .A1(n88), .A2(n107), .ZN(n666) );
  XNOR2_X1 U698 ( .A(n667), .B(n666), .ZN(n668) );
  AOI22_X1 U699 ( .A1(n668), .A2(n789), .B1(n745), .B2(f[9]), .ZN(n669) );
  INV_X1 U700 ( .A(n669), .ZN(n55) );
  INV_X1 U701 ( .A(n109), .ZN(n682) );
  NAND2_X1 U702 ( .A1(n682), .A2(n672), .ZN(n673) );
  XNOR2_X1 U703 ( .A(n674), .B(n673), .ZN(n675) );
  AOI22_X1 U704 ( .A1(n675), .A2(n789), .B1(n745), .B2(f[10]), .ZN(n788) );
  OR2_X1 U705 ( .A1(n677), .A2(n676), .ZN(n699) );
  NAND2_X1 U706 ( .A1(n699), .A2(n702), .ZN(n678) );
  XNOR2_X1 U707 ( .A(n679), .B(n678), .ZN(n680) );
  AOI22_X1 U708 ( .A1(n680), .A2(n789), .B1(n745), .B2(f[14]), .ZN(n681) );
  INV_X1 U709 ( .A(n681), .ZN(n50) );
  OAI21_X1 U710 ( .B1(n692), .B2(n109), .A(n672), .ZN(n687) );
  INV_X1 U711 ( .A(n683), .ZN(n685) );
  NAND2_X1 U712 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U713 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U714 ( .A1(n745), .A2(f[11]), .ZN(n689) );
  NAND2_X1 U715 ( .A1(n690), .A2(n689), .ZN(n53) );
  OAI21_X1 U716 ( .B1(n692), .B2(n145), .A(n691), .ZN(n695) );
  NAND2_X1 U717 ( .A1(n137), .A2(n118), .ZN(n694) );
  XNOR2_X1 U718 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U719 ( .A1(n745), .A2(f[12]), .ZN(n697) );
  NAND2_X1 U720 ( .A1(n698), .A2(n697), .ZN(n52) );
  INV_X1 U721 ( .A(n699), .ZN(n704) );
  NAND3_X1 U722 ( .A1(n700), .A2(n701), .A3(n699), .ZN(n703) );
  OAI211_X1 U723 ( .C1(n704), .C2(n705), .A(n703), .B(n702), .ZN(n710) );
  INV_X1 U724 ( .A(n706), .ZN(n708) );
  NAND2_X1 U725 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U726 ( .A(n710), .B(n709), .ZN(n711) );
  NAND2_X1 U727 ( .A1(n711), .A2(n789), .ZN(n713) );
  NAND2_X1 U728 ( .A1(n745), .A2(f[15]), .ZN(n712) );
  NAND2_X1 U729 ( .A1(n713), .A2(n712), .ZN(n49) );
  FA_X1 U730 ( .A(n716), .B(n715), .CI(n714), .CO(n729), .S(n557) );
  NOR2_X1 U731 ( .A1(n764), .A2(n142), .ZN(n717) );
  XOR2_X1 U732 ( .A(f[19]), .B(n717), .Z(n718) );
  XOR2_X1 U733 ( .A(f[18]), .B(n718), .Z(n727) );
  FA_X1 U734 ( .A(n720), .B(n765), .CI(n719), .CO(n725), .S(n716) );
  AOI21_X1 U735 ( .B1(n722), .B2(n128), .A(n764), .ZN(n723) );
  INV_X1 U736 ( .A(n723), .ZN(n724) );
  XOR2_X1 U737 ( .A(n725), .B(n724), .Z(n726) );
  XOR2_X1 U738 ( .A(n727), .B(n726), .Z(n728) );
  OR2_X1 U739 ( .A1(n729), .A2(n728), .ZN(n731) );
  NAND2_X1 U740 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U741 ( .A1(n731), .A2(n730), .ZN(n739) );
  INV_X1 U742 ( .A(n739), .ZN(n744) );
  NOR2_X1 U743 ( .A1(n732), .A2(n736), .ZN(n733) );
  NAND2_X1 U744 ( .A1(n734), .A2(n733), .ZN(n743) );
  OAI21_X1 U745 ( .B1(n737), .B2(n736), .A(n735), .ZN(n740) );
  INV_X1 U746 ( .A(n740), .ZN(n738) );
  NAND3_X1 U747 ( .A1(n743), .A2(n738), .A3(n744), .ZN(n742) );
  AOI21_X1 U748 ( .B1(n740), .B2(n739), .A(n530), .ZN(n741) );
  OAI211_X1 U749 ( .C1(n744), .C2(n743), .A(n742), .B(n741), .ZN(n747) );
  NAND2_X1 U750 ( .A1(n745), .A2(f[19]), .ZN(n746) );
  NAND2_X1 U751 ( .A1(n747), .A2(n746), .ZN(n45) );
  AOI22_X1 U752 ( .A1(n134), .A2(a[9]), .B1(n748), .B2(n752), .ZN(n774) );
  AOI22_X1 U753 ( .A1(n134), .A2(a[3]), .B1(n752), .B2(n96), .ZN(n775) );
  AOI22_X1 U754 ( .A1(n134), .A2(a[5]), .B1(n752), .B2(n115), .ZN(n776) );
  AOI22_X1 U755 ( .A1(n134), .A2(a[7]), .B1(n752), .B2(a_in[7]), .ZN(n777) );
  AOI22_X1 U756 ( .A1(n134), .A2(a[1]), .B1(n752), .B2(n102), .ZN(n778) );
endmodule

