
module part1_mac ( clk, reset, a, b, valid_in, f, valid_out );
  input [9:0] a;
  input [9:0] b;
  output [19:0] f;
  input clk, reset, valid_in;
  output valid_out;
  wire   enable_f, n47, n48, n49, n50, n51, n52, n53, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n77, n78, n79, n80, n82,
         n83, n86, \DP_OP_11J1_122_830/n421 , n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704;
  wire   [9:0] a_in;
  wire   [9:0] b_in;

  DFF_X1 \f_reg[19]  ( .D(n48), .CK(clk), .Q(f[19]), .QN(n686) );
  DFF_X1 \f_reg[18]  ( .D(n49), .CK(clk), .Q(f[18]) );
  DFF_X1 \f_reg[16]  ( .D(n51), .CK(clk), .Q(f[16]) );
  DFF_X1 \f_reg[14]  ( .D(n53), .CK(clk), .Q(f[14]) );
  DFF_X1 \f_reg[13]  ( .D(n668), .CK(clk), .Q(f[13]), .QN(n111) );
  DFF_X1 \f_reg[11]  ( .D(n56), .CK(clk), .Q(f[11]), .QN(n120) );
  DFF_X1 \a_in_reg[9]  ( .D(n77), .CK(clk), .Q(a_in[9]), .QN(n673) );
  DFF_X1 \a_in_reg[0]  ( .D(n86), .CK(clk), .Q(a_in[0]), .QN(n681) );
  DFF_X1 \b_in_reg[9]  ( .D(n68), .CK(clk), .Q(b_in[9]), .QN(n676) );
  DFF_X1 \f_reg[17]  ( .D(n50), .CK(clk), .Q(f[17]), .QN(n687) );
  DFF_X1 \b_in_reg[5]  ( .D(n700), .CK(clk), .Q(n690), .QN(
        \DP_OP_11J1_122_830/n421 ) );
  DFF_X1 \b_in_reg[1]  ( .D(n692), .CK(clk), .Q(n680), .QN(b_in[1]) );
  DFF_X1 \b_in_reg[8]  ( .D(n698), .CK(clk), .Q(n678), .QN(b_in[8]) );
  DFF_X1 \b_in_reg[3]  ( .D(n693), .CK(clk), .Q(n679), .QN(b_in[3]) );
  DFF_X1 \f_reg[15]  ( .D(n52), .CK(clk), .Q(f[15]), .QN(n688) );
  DFF_X1 \b_in_reg[7]  ( .D(n694), .CK(clk), .Q(n121), .QN(b_in[7]) );
  DFF_X1 \b_in_reg[2]  ( .D(n702), .CK(clk), .Q(n108), .QN(b_in[2]) );
  DFF_X1 enable_f_reg ( .D(n47), .CK(clk), .Q(enable_f), .QN(n691) );
  DFF_X1 \b_in_reg[6]  ( .D(n699), .CK(clk), .Q(n674), .QN(b_in[6]) );
  DFF_X1 valid_out_reg ( .D(n704), .CK(clk), .Q(valid_out) );
  DFF_X1 \f_reg[0]  ( .D(n67), .CK(clk), .Q(f[0]) );
  DFF_X1 \a_in_reg[8]  ( .D(n78), .CK(clk), .Q(a_in[8]) );
  DFF_X1 \a_in_reg[7]  ( .D(n79), .CK(clk), .Q(a_in[7]) );
  DFF_X1 \a_in_reg[6]  ( .D(n80), .CK(clk), .Q(a_in[6]) );
  DFF_X1 \a_in_reg[4]  ( .D(n82), .CK(clk), .Q(a_in[4]) );
  DFF_X1 \a_in_reg[3]  ( .D(n83), .CK(clk), .Q(a_in[3]) );
  DFF_X1 \f_reg[1]  ( .D(n66), .CK(clk), .Q(f[1]), .QN(n682) );
  DFF_X1 \f_reg[2]  ( .D(n65), .CK(clk), .Q(f[2]) );
  DFF_X1 \f_reg[3]  ( .D(n64), .CK(clk), .Q(f[3]), .QN(n685) );
  DFF_X1 \f_reg[4]  ( .D(n63), .CK(clk), .Q(f[4]) );
  DFF_X1 \f_reg[5]  ( .D(n62), .CK(clk), .Q(f[5]), .QN(n683) );
  DFF_X1 \f_reg[6]  ( .D(n61), .CK(clk), .Q(f[6]) );
  DFF_X1 \f_reg[7]  ( .D(n60), .CK(clk), .Q(f[7]) );
  DFF_X1 \f_reg[8]  ( .D(n59), .CK(clk), .Q(f[8]) );
  DFF_X1 \f_reg[9]  ( .D(n58), .CK(clk), .Q(f[9]), .QN(n684) );
  DFF_X1 \f_reg[10]  ( .D(n57), .CK(clk), .Q(f[10]) );
  DFF_X1 \a_in_reg[1]  ( .D(n697), .CK(clk), .Q(n675), .QN(a_in[1]) );
  DFF_X1 \a_in_reg[2]  ( .D(n696), .CK(clk), .Q(n677), .QN(a_in[2]) );
  DFFRS_X1 \f_reg[12]  ( .D(n55), .CK(clk), .RN(1'b1), .SN(1'b1), .Q(f[12]), 
        .QN(n113) );
  DFF_X1 \a_in_reg[5]  ( .D(n695), .CK(clk), .QN(a_in[5]) );
  DFF_X1 \b_in_reg[4]  ( .D(n701), .CK(clk), .Q(n104), .QN(b_in[4]) );
  DFF_X1 \b_in_reg[0]  ( .D(n703), .CK(clk), .Q(n689), .QN(b_in[0]) );
  OR2_X1 U91 ( .A1(b_in[0]), .A2(n680), .ZN(n437) );
  NOR2_X1 U92 ( .A1(n406), .A2(n405), .ZN(n602) );
  NAND2_X1 U93 ( .A1(n661), .A2(n660), .ZN(n88) );
  AOI21_X1 U94 ( .B1(n548), .B2(n550), .A(n194), .ZN(n554) );
  CLKBUF_X1 U95 ( .A(n520), .Z(n92) );
  OR2_X1 U96 ( .A1(n527), .A2(n531), .ZN(n232) );
  CLKBUF_X1 U97 ( .A(n337), .Z(n107) );
  CLKBUF_X1 U98 ( .A(n272), .Z(n96) );
  AND2_X1 U99 ( .A1(n374), .A2(f[3]), .ZN(n393) );
  BUF_X1 U100 ( .A(n416), .Z(n89) );
  INV_X1 U101 ( .A(n121), .ZN(n90) );
  BUF_X1 U102 ( .A(n284), .Z(n91) );
  AOI21_X1 U103 ( .B1(n99), .B2(n536), .A(n535), .ZN(n657) );
  NOR2_X1 U104 ( .A1(n553), .A2(n232), .ZN(n93) );
  INV_X1 U105 ( .A(n163), .ZN(n94) );
  BUF_X1 U106 ( .A(n416), .Z(n95) );
  AND2_X1 U107 ( .A1(n322), .A2(n321), .ZN(n97) );
  BUF_X1 U108 ( .A(n679), .Z(n98) );
  NAND2_X1 U109 ( .A1(n456), .A2(n616), .ZN(n99) );
  BUF_X1 U110 ( .A(n586), .Z(n100) );
  BUF_X1 U111 ( .A(n653), .Z(n101) );
  NOR2_X1 U112 ( .A1(n490), .A2(n489), .ZN(n102) );
  NOR2_X1 U113 ( .A1(n490), .A2(n489), .ZN(n103) );
  INV_X1 U114 ( .A(n353), .ZN(n355) );
  XNOR2_X1 U115 ( .A(n104), .B(\DP_OP_11J1_122_830/n421 ), .ZN(n135) );
  BUF_X1 U116 ( .A(n657), .Z(n105) );
  BUF_X1 U117 ( .A(n344), .Z(n106) );
  XNOR2_X1 U118 ( .A(n108), .B(b_in[3]), .ZN(n136) );
  XNOR2_X1 U119 ( .A(n339), .B(n338), .ZN(n109) );
  XOR2_X1 U120 ( .A(n98), .B(a_in[8]), .Z(n234) );
  XNOR2_X1 U121 ( .A(b_in[4]), .B(n679), .ZN(n353) );
  BUF_X1 U122 ( .A(n655), .Z(n110) );
  NOR2_X1 U123 ( .A1(n349), .A2(n348), .ZN(n655) );
  OAI22_X1 U124 ( .A1(n371), .A2(n414), .B1(n416), .B2(n370), .ZN(n401) );
  XNOR2_X1 U125 ( .A(f[11]), .B(f[12]), .ZN(n166) );
  AND2_X1 U126 ( .A1(n417), .A2(f[5]), .ZN(n443) );
  INV_X1 U127 ( .A(n401), .ZN(n398) );
  OR2_X1 U128 ( .A1(n263), .A2(f[10]), .ZN(n252) );
  INV_X1 U129 ( .A(n180), .ZN(n150) );
  XNOR2_X1 U130 ( .A(n385), .B(n682), .ZN(n576) );
  NAND2_X1 U131 ( .A1(n243), .A2(n242), .ZN(n282) );
  XNOR2_X1 U132 ( .A(n308), .B(n307), .ZN(n459) );
  XNOR2_X1 U133 ( .A(n306), .B(n305), .ZN(n308) );
  CLKBUF_X1 U134 ( .A(n463), .Z(n464) );
  INV_X1 U135 ( .A(n484), .ZN(n480) );
  INV_X1 U136 ( .A(n483), .ZN(n479) );
  INV_X1 U137 ( .A(n428), .ZN(n424) );
  INV_X1 U138 ( .A(n429), .ZN(n425) );
  INV_X1 U139 ( .A(n393), .ZN(n366) );
  INV_X1 U140 ( .A(n394), .ZN(n365) );
  XNOR2_X1 U141 ( .A(n329), .B(n328), .ZN(n342) );
  XNOR2_X1 U142 ( .A(n327), .B(n326), .ZN(n329) );
  NAND2_X1 U143 ( .A1(n176), .A2(n175), .ZN(n338) );
  NAND2_X1 U144 ( .A1(n327), .A2(n326), .ZN(n175) );
  NAND2_X1 U145 ( .A1(n486), .A2(n485), .ZN(n487) );
  NAND2_X1 U146 ( .A1(n484), .A2(n483), .ZN(n485) );
  NAND2_X1 U147 ( .A1(n482), .A2(n481), .ZN(n486) );
  NAND2_X1 U148 ( .A1(n480), .A2(n479), .ZN(n481) );
  NOR2_X1 U149 ( .A1(n488), .A2(n487), .ZN(n628) );
  NAND2_X1 U150 ( .A1(n452), .A2(n451), .ZN(n454) );
  NAND2_X1 U151 ( .A1(n448), .A2(n447), .ZN(n452) );
  NAND2_X1 U152 ( .A1(n431), .A2(n430), .ZN(n432) );
  NAND2_X1 U153 ( .A1(n429), .A2(n428), .ZN(n430) );
  NAND2_X1 U154 ( .A1(n427), .A2(n426), .ZN(n431) );
  NAND2_X1 U155 ( .A1(n425), .A2(n424), .ZN(n426) );
  NAND2_X1 U156 ( .A1(n369), .A2(n368), .ZN(n407) );
  NAND2_X1 U157 ( .A1(n393), .A2(n394), .ZN(n368) );
  NAND2_X1 U158 ( .A1(n396), .A2(n367), .ZN(n369) );
  NAND2_X1 U159 ( .A1(n366), .A2(n365), .ZN(n367) );
  NAND2_X1 U160 ( .A1(n404), .A2(n403), .ZN(n405) );
  NAND2_X1 U161 ( .A1(n400), .A2(n399), .ZN(n404) );
  NAND2_X1 U162 ( .A1(n398), .A2(n397), .ZN(n400) );
  NAND2_X1 U163 ( .A1(n380), .A2(n379), .ZN(n391) );
  NAND2_X1 U164 ( .A1(n382), .A2(f[2]), .ZN(n379) );
  AND2_X1 U165 ( .A1(n392), .A2(n391), .ZN(n582) );
  AND2_X1 U166 ( .A1(n385), .A2(f[1]), .ZN(n389) );
  NAND2_X1 U167 ( .A1(n314), .A2(n313), .ZN(n287) );
  NAND2_X1 U168 ( .A1(n333), .A2(n332), .ZN(n335) );
  NAND2_X1 U169 ( .A1(n182), .A2(n181), .ZN(n229) );
  NAND2_X1 U170 ( .A1(n338), .A2(n336), .ZN(n181) );
  OAI21_X1 U171 ( .B1(n336), .B2(n338), .A(n107), .ZN(n182) );
  OAI21_X1 U172 ( .B1(n150), .B2(n149), .A(n148), .ZN(n191) );
  OR2_X1 U173 ( .A1(n529), .A2(n531), .ZN(n222) );
  INV_X1 U174 ( .A(n220), .ZN(n221) );
  OAI21_X1 U175 ( .B1(n528), .B2(n531), .A(n532), .ZN(n220) );
  INV_X1 U176 ( .A(n582), .ZN(n583) );
  OAI22_X1 U177 ( .A1(n576), .A2(n122), .B1(n575), .B2(n388), .ZN(n593) );
  INV_X1 U178 ( .A(n578), .ZN(n388) );
  NAND2_X1 U179 ( .A1(n576), .A2(n575), .ZN(n577) );
  AND2_X1 U180 ( .A1(valid_in), .A2(n563), .ZN(n671) );
  OR2_X1 U181 ( .A1(n501), .A2(n503), .ZN(n506) );
  AND2_X1 U182 ( .A1(n662), .A2(f[13]), .ZN(n112) );
  NOR2_X1 U183 ( .A1(n553), .A2(n527), .ZN(n114) );
  NAND2_X1 U184 ( .A1(n609), .A2(n596), .ZN(n115) );
  AND2_X1 U185 ( .A1(enable_f), .A2(n563), .ZN(n704) );
  NAND2_X1 U186 ( .A1(n559), .A2(n558), .ZN(n116) );
  NAND2_X1 U187 ( .A1(n231), .A2(n532), .ZN(n117) );
  NAND2_X1 U188 ( .A1(n544), .A2(n543), .ZN(n118) );
  NAND2_X1 U189 ( .A1(n550), .A2(n549), .ZN(n119) );
  AND2_X1 U190 ( .A1(n575), .A2(n388), .ZN(n122) );
  AND2_X1 U191 ( .A1(n88), .A2(n704), .ZN(n123) );
  OR2_X1 U192 ( .A1(n576), .A2(n575), .ZN(n124) );
  OR2_X1 U193 ( .A1(n656), .A2(n110), .ZN(n125) );
  NOR2_X1 U194 ( .A1(n553), .A2(n232), .ZN(n126) );
  NAND2_X1 U195 ( .A1(n662), .A2(f[18]), .ZN(n127) );
  NAND2_X1 U196 ( .A1(n662), .A2(f[17]), .ZN(n128) );
  NAND2_X1 U197 ( .A1(n662), .A2(f[15]), .ZN(n129) );
  NAND2_X1 U198 ( .A1(n662), .A2(f[16]), .ZN(n130) );
  NAND2_X1 U199 ( .A1(n662), .A2(f[19]), .ZN(n131) );
  OR2_X1 U200 ( .A1(n433), .A2(n432), .ZN(n615) );
  OR2_X1 U201 ( .A1(n88), .A2(n546), .ZN(n132) );
  INV_X1 U203 ( .A(reset), .ZN(n563) );
  XOR2_X1 U204 ( .A(n90), .B(b_in[6]), .Z(n133) );
  XNOR2_X1 U205 ( .A(n690), .B(n674), .ZN(n170) );
  NAND2_X2 U206 ( .A1(n133), .A2(n170), .ZN(n296) );
  BUF_X2 U207 ( .A(b_in[7]), .Z(n292) );
  XNOR2_X1 U208 ( .A(n292), .B(a_in[5]), .ZN(n171) );
  XNOR2_X1 U209 ( .A(n292), .B(a_in[6]), .ZN(n147) );
  OAI22_X1 U210 ( .A1(n296), .A2(n171), .B1(n294), .B2(n147), .ZN(n325) );
  XNOR2_X1 U211 ( .A(b_in[3]), .B(b_in[4]), .ZN(n134) );
  NAND2_X2 U212 ( .A1(n135), .A2(n134), .ZN(n412) );
  INV_X2 U213 ( .A(n690), .ZN(n669) );
  XNOR2_X1 U214 ( .A(n669), .B(a_in[7]), .ZN(n172) );
  XNOR2_X1 U215 ( .A(n669), .B(a_in[8]), .ZN(n157) );
  OAI22_X1 U216 ( .A1(n412), .A2(n172), .B1(n355), .B2(n157), .ZN(n324) );
  XNOR2_X1 U217 ( .A(n98), .B(n673), .ZN(n161) );
  INV_X1 U218 ( .A(n161), .ZN(n139) );
  XNOR2_X1 U219 ( .A(b_in[1]), .B(b_in[2]), .ZN(n137) );
  BUF_X2 U220 ( .A(n137), .Z(n414) );
  NAND2_X2 U221 ( .A1(n137), .A2(n136), .ZN(n416) );
  NAND2_X1 U222 ( .A1(n414), .A2(n416), .ZN(n138) );
  NAND2_X1 U223 ( .A1(n139), .A2(n138), .ZN(n323) );
  NAND2_X1 U224 ( .A1(n120), .A2(n113), .ZN(n140) );
  XNOR2_X1 U225 ( .A(b_in[7]), .B(b_in[8]), .ZN(n142) );
  XNOR2_X1 U226 ( .A(b_in[9]), .B(n678), .ZN(n141) );
  NAND2_X2 U227 ( .A1(n142), .A2(n141), .ZN(n249) );
  INV_X1 U228 ( .A(n249), .ZN(n163) );
  NAND2_X1 U229 ( .A1(n140), .A2(n163), .ZN(n146) );
  BUF_X2 U230 ( .A(b_in[9]), .Z(n650) );
  XNOR2_X1 U231 ( .A(n650), .B(a_in[3]), .ZN(n160) );
  INV_X1 U232 ( .A(n160), .ZN(n162) );
  XNOR2_X1 U233 ( .A(n650), .B(a_in[4]), .ZN(n155) );
  BUF_X1 U234 ( .A(n142), .Z(n247) );
  OR2_X1 U235 ( .A1(n155), .A2(n247), .ZN(n164) );
  INV_X1 U236 ( .A(n164), .ZN(n143) );
  NAND2_X1 U237 ( .A1(n143), .A2(n140), .ZN(n145) );
  NAND2_X1 U238 ( .A1(f[11]), .A2(f[12]), .ZN(n144) );
  OAI211_X1 U239 ( .C1(n146), .C2(n160), .A(n145), .B(n144), .ZN(n178) );
  XNOR2_X1 U240 ( .A(n292), .B(a_in[7]), .ZN(n152) );
  OAI22_X1 U241 ( .A1(n296), .A2(n147), .B1(n294), .B2(n152), .ZN(n177) );
  NOR2_X1 U242 ( .A1(n178), .A2(n177), .ZN(n149) );
  NAND2_X1 U243 ( .A1(n178), .A2(n177), .ZN(n148) );
  XOR2_X1 U244 ( .A(n676), .B(a_in[5]), .Z(n154) );
  INV_X1 U245 ( .A(n237), .ZN(n269) );
  INV_X1 U246 ( .A(n676), .ZN(n246) );
  XNOR2_X1 U247 ( .A(n246), .B(a_in[6]), .ZN(n183) );
  OAI22_X1 U248 ( .A1(n94), .A2(n154), .B1(n237), .B2(n183), .ZN(n185) );
  INV_X1 U249 ( .A(n353), .ZN(n410) );
  XNOR2_X1 U250 ( .A(n669), .B(a_in[9]), .ZN(n156) );
  AOI21_X1 U251 ( .B1(n412), .B2(n410), .A(n156), .ZN(n151) );
  INV_X1 U252 ( .A(n151), .ZN(n188) );
  XNOR2_X1 U253 ( .A(n292), .B(a_in[8]), .ZN(n184) );
  OAI22_X1 U254 ( .A1(n296), .A2(n152), .B1(n294), .B2(n184), .ZN(n187) );
  XNOR2_X1 U255 ( .A(b_in[7]), .B(b_in[8]), .ZN(n153) );
  BUF_X2 U256 ( .A(n153), .Z(n237) );
  OAI22_X1 U257 ( .A1(n249), .A2(n155), .B1(n237), .B2(n154), .ZN(n159) );
  OAI22_X1 U258 ( .A1(n412), .A2(n157), .B1(n410), .B2(n156), .ZN(n158) );
  FA_X1 U259 ( .A(n159), .B(n111), .CI(n158), .CO(n186), .S(n336) );
  XNOR2_X1 U260 ( .A(n676), .B(n677), .ZN(n173) );
  OAI22_X1 U261 ( .A1(n249), .A2(n173), .B1(n237), .B2(n160), .ZN(n256) );
  BUF_X2 U262 ( .A(b_in[3]), .Z(n652) );
  OAI22_X1 U263 ( .A1(n416), .A2(n234), .B1(n414), .B2(n161), .ZN(n255) );
  INV_X1 U264 ( .A(n327), .ZN(n169) );
  NAND2_X1 U265 ( .A1(n163), .A2(n162), .ZN(n165) );
  NAND2_X1 U266 ( .A1(n165), .A2(n164), .ZN(n167) );
  XNOR2_X1 U267 ( .A(n167), .B(n166), .ZN(n326) );
  INV_X1 U268 ( .A(n326), .ZN(n168) );
  NAND2_X1 U269 ( .A1(n169), .A2(n168), .ZN(n174) );
  XNOR2_X1 U270 ( .A(n292), .B(a_in[4]), .ZN(n261) );
  BUF_X2 U271 ( .A(n170), .Z(n294) );
  OAI22_X1 U272 ( .A1(n296), .A2(n261), .B1(n294), .B2(n171), .ZN(n254) );
  XNOR2_X1 U273 ( .A(\DP_OP_11J1_122_830/n421 ), .B(a_in[6]), .ZN(n235) );
  OAI22_X1 U274 ( .A1(n412), .A2(n235), .B1(n355), .B2(n172), .ZN(n253) );
  XNOR2_X1 U275 ( .A(n676), .B(n675), .ZN(n236) );
  OAI22_X1 U276 ( .A1(n249), .A2(n236), .B1(n247), .B2(n173), .ZN(n263) );
  NAND2_X1 U277 ( .A1(n174), .A2(n328), .ZN(n176) );
  XNOR2_X1 U278 ( .A(n178), .B(n177), .ZN(n179) );
  XNOR2_X1 U279 ( .A(n179), .B(n180), .ZN(n337) );
  NAND2_X1 U280 ( .A1(n230), .A2(n229), .ZN(n643) );
  INV_X1 U281 ( .A(n643), .ZN(n548) );
  XNOR2_X1 U282 ( .A(n650), .B(a_in[7]), .ZN(n199) );
  OAI22_X1 U283 ( .A1(n94), .A2(n183), .B1(n237), .B2(n199), .ZN(n196) );
  XNOR2_X1 U284 ( .A(n292), .B(a_in[9]), .ZN(n197) );
  OAI22_X1 U285 ( .A1(n296), .A2(n184), .B1(n294), .B2(n197), .ZN(n195) );
  FA_X1 U286 ( .A(f[13]), .B(f[14]), .CI(n185), .CO(n201), .S(n190) );
  FA_X1 U287 ( .A(n188), .B(n187), .CI(n186), .CO(n200), .S(n189) );
  FA_X1 U288 ( .A(n191), .B(n190), .CI(n189), .CO(n192), .S(n230) );
  OR2_X1 U289 ( .A1(n193), .A2(n192), .ZN(n550) );
  NAND2_X1 U290 ( .A1(n193), .A2(n192), .ZN(n549) );
  INV_X1 U291 ( .A(n549), .ZN(n194) );
  FA_X1 U292 ( .A(n196), .B(n688), .CI(n195), .CO(n207), .S(n202) );
  AOI21_X1 U293 ( .B1(n294), .B2(n296), .A(n197), .ZN(n198) );
  INV_X1 U294 ( .A(n198), .ZN(n206) );
  XNOR2_X1 U295 ( .A(n650), .B(a_in[8]), .ZN(n203) );
  OAI22_X1 U296 ( .A1(n249), .A2(n199), .B1(n237), .B2(n203), .ZN(n204) );
  FA_X1 U297 ( .A(n202), .B(n201), .CI(n200), .CO(n212), .S(n193) );
  NOR2_X1 U298 ( .A1(n213), .A2(n212), .ZN(n540) );
  XNOR2_X1 U299 ( .A(n246), .B(a_in[9]), .ZN(n210) );
  OAI22_X1 U300 ( .A1(n94), .A2(n203), .B1(n153), .B2(n210), .ZN(n209) );
  FA_X1 U301 ( .A(f[15]), .B(f[16]), .CI(n204), .CO(n208), .S(n205) );
  FA_X1 U302 ( .A(n207), .B(n206), .CI(n205), .CO(n214), .S(n213) );
  OR2_X1 U303 ( .A1(n215), .A2(n214), .ZN(n544) );
  INV_X1 U304 ( .A(n544), .ZN(n216) );
  OR2_X1 U305 ( .A1(n540), .A2(n216), .ZN(n529) );
  FA_X1 U306 ( .A(n209), .B(n687), .CI(n208), .CO(n219), .S(n215) );
  AOI21_X1 U307 ( .B1(n237), .B2(n94), .A(n210), .ZN(n211) );
  INV_X1 U308 ( .A(n211), .ZN(n223) );
  NOR2_X1 U309 ( .A1(n219), .A2(n218), .ZN(n531) );
  NAND2_X1 U310 ( .A1(n213), .A2(n212), .ZN(n558) );
  NAND2_X1 U311 ( .A1(n215), .A2(n214), .ZN(n543) );
  OAI21_X1 U312 ( .B1(n558), .B2(n216), .A(n543), .ZN(n217) );
  INV_X1 U313 ( .A(n217), .ZN(n528) );
  NAND2_X1 U314 ( .A1(n219), .A2(n218), .ZN(n532) );
  OAI21_X1 U315 ( .B1(n554), .B2(n222), .A(n221), .ZN(n499) );
  INV_X1 U316 ( .A(n499), .ZN(n227) );
  FA_X1 U317 ( .A(f[17]), .B(f[18]), .CI(n223), .CO(n224), .S(n218) );
  OR2_X1 U318 ( .A1(n224), .A2(n686), .ZN(n226) );
  NAND2_X1 U319 ( .A1(n224), .A2(n686), .ZN(n225) );
  AND2_X1 U320 ( .A1(n226), .A2(n225), .ZN(n498) );
  INV_X1 U321 ( .A(n498), .ZN(n503) );
  OAI21_X1 U322 ( .B1(n227), .B2(n503), .A(n704), .ZN(n228) );
  INV_X1 U323 ( .A(n228), .ZN(n508) );
  OR2_X1 U324 ( .A1(n230), .A2(n229), .ZN(n644) );
  NAND2_X1 U325 ( .A1(n644), .A2(n550), .ZN(n553) );
  INV_X1 U326 ( .A(n540), .ZN(n559) );
  NAND2_X1 U327 ( .A1(n559), .A2(n544), .ZN(n527) );
  INV_X1 U328 ( .A(n531), .ZN(n231) );
  INV_X1 U329 ( .A(n680), .ZN(n362) );
  XNOR2_X1 U330 ( .A(n362), .B(a_in[9]), .ZN(n239) );
  AOI21_X1 U331 ( .B1(n437), .B2(n689), .A(n239), .ZN(n233) );
  INV_X1 U332 ( .A(n233), .ZN(n259) );
  XNOR2_X1 U333 ( .A(n652), .B(a_in[7]), .ZN(n245) );
  OAI22_X1 U334 ( .A1(n416), .A2(n245), .B1(n414), .B2(n234), .ZN(n258) );
  XNOR2_X1 U335 ( .A(n669), .B(a_in[5]), .ZN(n244) );
  OAI22_X1 U336 ( .A1(n412), .A2(n244), .B1(n410), .B2(n235), .ZN(n257) );
  XNOR2_X1 U337 ( .A(n292), .B(a_in[2]), .ZN(n266) );
  XNOR2_X1 U338 ( .A(n292), .B(a_in[3]), .ZN(n262) );
  OAI22_X1 U339 ( .A1(n296), .A2(n266), .B1(n294), .B2(n262), .ZN(n273) );
  XNOR2_X1 U340 ( .A(n246), .B(a_in[0]), .ZN(n238) );
  OAI22_X1 U341 ( .A1(n249), .A2(n238), .B1(n237), .B2(n236), .ZN(n272) );
  BUF_X2 U342 ( .A(b_in[1]), .Z(n649) );
  XNOR2_X1 U343 ( .A(n649), .B(a_in[8]), .ZN(n270) );
  OR2_X1 U344 ( .A1(n239), .A2(n689), .ZN(n240) );
  OAI21_X1 U345 ( .B1(n270), .B2(n437), .A(n240), .ZN(n271) );
  OR2_X1 U346 ( .A1(n272), .A2(n271), .ZN(n241) );
  NAND2_X1 U347 ( .A1(n273), .A2(n241), .ZN(n243) );
  NAND2_X1 U348 ( .A1(n96), .A2(n271), .ZN(n242) );
  XNOR2_X1 U349 ( .A(n669), .B(a_in[4]), .ZN(n268) );
  OAI22_X1 U350 ( .A1(n412), .A2(n268), .B1(n410), .B2(n244), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n652), .B(a_in[6]), .ZN(n267) );
  OAI22_X1 U352 ( .A1(n89), .A2(n267), .B1(n414), .B2(n245), .ZN(n302) );
  OR2_X1 U353 ( .A1(a_in[0]), .A2(n676), .ZN(n248) );
  OAI22_X1 U354 ( .A1(n249), .A2(n676), .B1(n248), .B2(n247), .ZN(n260) );
  XNOR2_X1 U355 ( .A(n260), .B(n684), .ZN(n301) );
  OAI21_X1 U356 ( .B1(n284), .B2(n282), .A(n283), .ZN(n251) );
  NAND2_X1 U357 ( .A1(n284), .A2(n282), .ZN(n250) );
  NAND2_X1 U358 ( .A1(n251), .A2(n250), .ZN(n333) );
  FA_X1 U359 ( .A(n254), .B(n253), .CI(n252), .CO(n328), .S(n332) );
  XNOR2_X1 U360 ( .A(n333), .B(n332), .ZN(n265) );
  FA_X1 U361 ( .A(n120), .B(n255), .CI(n256), .CO(n327), .S(n320) );
  FA_X1 U362 ( .A(n259), .B(n258), .CI(n257), .CO(n319), .S(n284) );
  XNOR2_X1 U363 ( .A(n320), .B(n319), .ZN(n264) );
  AND2_X1 U364 ( .A1(n260), .A2(f[9]), .ZN(n279) );
  OAI22_X1 U365 ( .A1(n296), .A2(n262), .B1(n294), .B2(n261), .ZN(n278) );
  XNOR2_X1 U366 ( .A(n263), .B(f[10]), .ZN(n277) );
  XNOR2_X1 U367 ( .A(n264), .B(n318), .ZN(n331) );
  XNOR2_X1 U368 ( .A(n265), .B(n331), .ZN(n494) );
  XNOR2_X1 U369 ( .A(n292), .B(a_in[1]), .ZN(n293) );
  OAI22_X1 U370 ( .A1(n296), .A2(n293), .B1(n294), .B2(n266), .ZN(n471) );
  XNOR2_X1 U371 ( .A(n652), .B(a_in[5]), .ZN(n291) );
  OAI22_X1 U372 ( .A1(n416), .A2(n291), .B1(n414), .B2(n267), .ZN(n470) );
  XNOR2_X1 U373 ( .A(\DP_OP_11J1_122_830/n421 ), .B(a_in[3]), .ZN(n290) );
  OAI22_X1 U374 ( .A1(n412), .A2(n290), .B1(n355), .B2(n268), .ZN(n469) );
  AND2_X1 U375 ( .A1(a_in[0]), .A2(n269), .ZN(n298) );
  XNOR2_X1 U376 ( .A(n649), .B(a_in[7]), .ZN(n435) );
  OAI22_X1 U377 ( .A1(n437), .A2(n435), .B1(n270), .B2(n689), .ZN(n297) );
  XNOR2_X1 U378 ( .A(n272), .B(n271), .ZN(n274) );
  XNOR2_X1 U379 ( .A(n274), .B(n273), .ZN(n307) );
  OAI21_X1 U380 ( .B1(n306), .B2(n305), .A(n307), .ZN(n276) );
  NAND2_X1 U381 ( .A1(n306), .A2(n305), .ZN(n275) );
  NAND2_X1 U382 ( .A1(n276), .A2(n275), .ZN(n314) );
  INV_X1 U383 ( .A(n314), .ZN(n281) );
  FA_X1 U384 ( .A(n279), .B(n278), .CI(n277), .CO(n318), .S(n313) );
  INV_X1 U385 ( .A(n313), .ZN(n280) );
  NAND2_X1 U386 ( .A1(n281), .A2(n280), .ZN(n286) );
  XNOR2_X1 U387 ( .A(n283), .B(n282), .ZN(n285) );
  XNOR2_X1 U388 ( .A(n285), .B(n91), .ZN(n315) );
  NAND2_X1 U389 ( .A1(n286), .A2(n315), .ZN(n288) );
  NAND2_X1 U390 ( .A1(n288), .A2(n287), .ZN(n493) );
  NOR2_X1 U391 ( .A1(n494), .A2(n493), .ZN(n317) );
  NAND2_X1 U392 ( .A1(n292), .A2(n681), .ZN(n289) );
  OAI22_X1 U393 ( .A1(n294), .A2(n289), .B1(n296), .B2(n121), .ZN(n442) );
  XNOR2_X1 U394 ( .A(n669), .B(a_in[2]), .ZN(n409) );
  OAI22_X1 U395 ( .A1(n412), .A2(n409), .B1(n355), .B2(n290), .ZN(n441) );
  XNOR2_X1 U396 ( .A(n652), .B(a_in[4]), .ZN(n413) );
  OAI22_X1 U397 ( .A1(n416), .A2(n413), .B1(n414), .B2(n291), .ZN(n440) );
  XNOR2_X1 U398 ( .A(n292), .B(a_in[0]), .ZN(n295) );
  OAI22_X1 U399 ( .A1(n296), .A2(n295), .B1(n294), .B2(n293), .ZN(n434) );
  FA_X1 U400 ( .A(n298), .B(f[8]), .CI(n297), .CO(n305), .S(n463) );
  OAI21_X1 U401 ( .B1(n462), .B2(n461), .A(n463), .ZN(n300) );
  NAND2_X1 U402 ( .A1(n462), .A2(n461), .ZN(n299) );
  NAND2_X1 U403 ( .A1(n300), .A2(n299), .ZN(n457) );
  INV_X1 U404 ( .A(n457), .ZN(n304) );
  FA_X1 U405 ( .A(n303), .B(n302), .CI(n301), .CO(n283), .S(n458) );
  INV_X1 U406 ( .A(n458), .ZN(n310) );
  NAND2_X1 U407 ( .A1(n304), .A2(n310), .ZN(n309) );
  NAND2_X1 U408 ( .A1(n309), .A2(n459), .ZN(n312) );
  NAND2_X1 U409 ( .A1(n457), .A2(n458), .ZN(n311) );
  NAND2_X1 U410 ( .A1(n312), .A2(n311), .ZN(n492) );
  XNOR2_X1 U411 ( .A(n314), .B(n313), .ZN(n316) );
  XNOR2_X1 U412 ( .A(n316), .B(n315), .ZN(n491) );
  NAND2_X1 U413 ( .A1(n492), .A2(n491), .ZN(n637) );
  NAND2_X1 U414 ( .A1(n494), .A2(n493), .ZN(n521) );
  OAI21_X1 U415 ( .B1(n317), .B2(n637), .A(n521), .ZN(n510) );
  OAI21_X1 U416 ( .B1(n320), .B2(n319), .A(n318), .ZN(n322) );
  NAND2_X1 U417 ( .A1(n320), .A2(n319), .ZN(n321) );
  NAND2_X1 U418 ( .A1(n322), .A2(n321), .ZN(n344) );
  FA_X1 U419 ( .A(n325), .B(n324), .CI(n323), .CO(n180), .S(n343) );
  XNOR2_X1 U420 ( .A(n344), .B(n343), .ZN(n330) );
  XNOR2_X1 U421 ( .A(n330), .B(n342), .ZN(n349) );
  OAI21_X1 U422 ( .B1(n333), .B2(n332), .A(n331), .ZN(n334) );
  NAND2_X1 U423 ( .A1(n334), .A2(n335), .ZN(n348) );
  XNOR2_X1 U424 ( .A(n337), .B(n336), .ZN(n339) );
  XNOR2_X1 U425 ( .A(n339), .B(n338), .ZN(n659) );
  INV_X1 U426 ( .A(n343), .ZN(n340) );
  NAND2_X1 U427 ( .A1(n97), .A2(n340), .ZN(n341) );
  NAND2_X1 U428 ( .A1(n341), .A2(n342), .ZN(n346) );
  NAND2_X1 U429 ( .A1(n106), .A2(n343), .ZN(n345) );
  NAND2_X1 U430 ( .A1(n346), .A2(n345), .ZN(n658) );
  NOR2_X1 U431 ( .A1(n109), .A2(n658), .ZN(n347) );
  NOR2_X1 U432 ( .A1(n347), .A2(n655), .ZN(n495) );
  NOR2_X1 U433 ( .A1(n659), .A2(n658), .ZN(n350) );
  NAND2_X1 U434 ( .A1(n349), .A2(n348), .ZN(n653) );
  NAND2_X1 U435 ( .A1(n659), .A2(n658), .ZN(n660) );
  OAI21_X1 U436 ( .B1(n350), .B2(n653), .A(n660), .ZN(n351) );
  AOI21_X1 U437 ( .B1(n510), .B2(n495), .A(n351), .ZN(n537) );
  INV_X1 U438 ( .A(n537), .ZN(n352) );
  NAND2_X1 U439 ( .A1(n93), .A2(n352), .ZN(n501) );
  AND2_X1 U440 ( .A1(a_in[0]), .A2(n353), .ZN(n361) );
  XNOR2_X1 U441 ( .A(n649), .B(a_in[3]), .ZN(n363) );
  XNOR2_X1 U442 ( .A(n649), .B(a_in[4]), .ZN(n358) );
  OAI22_X1 U443 ( .A1(n437), .A2(n363), .B1(n358), .B2(n689), .ZN(n360) );
  XNOR2_X1 U444 ( .A(n669), .B(a_in[0]), .ZN(n354) );
  XNOR2_X1 U445 ( .A(n669), .B(a_in[1]), .ZN(n411) );
  OAI22_X1 U446 ( .A1(n412), .A2(n354), .B1(n410), .B2(n411), .ZN(n417) );
  XNOR2_X1 U447 ( .A(n417), .B(n683), .ZN(n428) );
  XNOR2_X1 U448 ( .A(n429), .B(n428), .ZN(n359) );
  INV_X1 U449 ( .A(n669), .ZN(n357) );
  OR2_X1 U450 ( .A1(a_in[0]), .A2(n357), .ZN(n356) );
  OAI22_X1 U451 ( .A1(n412), .A2(n357), .B1(n356), .B2(n355), .ZN(n422) );
  XNOR2_X1 U452 ( .A(n649), .B(a_in[5]), .ZN(n418) );
  OAI22_X1 U453 ( .A1(n437), .A2(n358), .B1(n418), .B2(n689), .ZN(n421) );
  XNOR2_X1 U454 ( .A(n652), .B(a_in[2]), .ZN(n364) );
  XNOR2_X1 U455 ( .A(n652), .B(a_in[3]), .ZN(n415) );
  OAI22_X1 U456 ( .A1(n95), .A2(n364), .B1(n414), .B2(n415), .ZN(n420) );
  XNOR2_X1 U457 ( .A(n359), .B(n427), .ZN(n408) );
  FA_X1 U458 ( .A(n361), .B(f[4]), .CI(n360), .CO(n429), .S(n396) );
  XNOR2_X1 U459 ( .A(n362), .B(a_in[2]), .ZN(n377) );
  OAI22_X1 U460 ( .A1(n363), .A2(n689), .B1(n437), .B2(n377), .ZN(n374) );
  XNOR2_X1 U461 ( .A(n652), .B(a_in[1]), .ZN(n372) );
  OAI22_X1 U462 ( .A1(n89), .A2(n372), .B1(n414), .B2(n364), .ZN(n394) );
  NAND2_X1 U463 ( .A1(n408), .A2(n407), .ZN(n596) );
  NAND2_X1 U464 ( .A1(n652), .A2(n681), .ZN(n371) );
  INV_X1 U465 ( .A(n652), .ZN(n370) );
  XNOR2_X1 U466 ( .A(n652), .B(a_in[0]), .ZN(n373) );
  OAI22_X1 U467 ( .A1(n416), .A2(n373), .B1(n414), .B2(n372), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n401), .B(n402), .ZN(n375) );
  XNOR2_X1 U469 ( .A(n374), .B(n685), .ZN(n399) );
  XNOR2_X1 U470 ( .A(n375), .B(n399), .ZN(n392) );
  INV_X1 U471 ( .A(n414), .ZN(n376) );
  AND2_X1 U472 ( .A1(a_in[0]), .A2(n376), .ZN(n382) );
  XNOR2_X1 U473 ( .A(n649), .B(a_in[1]), .ZN(n384) );
  OR2_X1 U474 ( .A1(n377), .A2(n689), .ZN(n378) );
  OAI21_X1 U475 ( .B1(n384), .B2(n437), .A(n378), .ZN(n381) );
  OAI21_X1 U476 ( .B1(n382), .B2(f[2]), .A(n381), .ZN(n380) );
  OR2_X1 U477 ( .A1(n392), .A2(n391), .ZN(n584) );
  XNOR2_X1 U478 ( .A(n381), .B(f[2]), .ZN(n383) );
  XNOR2_X1 U479 ( .A(n383), .B(n382), .ZN(n390) );
  OAI22_X1 U480 ( .A1(n384), .A2(n689), .B1(n437), .B2(a_in[0]), .ZN(n385) );
  NOR2_X1 U481 ( .A1(n390), .A2(n389), .ZN(n589) );
  INV_X1 U482 ( .A(n649), .ZN(n386) );
  OR2_X1 U483 ( .A1(a_in[0]), .A2(n386), .ZN(n387) );
  NAND2_X1 U484 ( .A1(n387), .A2(n437), .ZN(n575) );
  AND2_X1 U485 ( .A1(a_in[0]), .A2(b_in[0]), .ZN(n564) );
  NAND2_X1 U486 ( .A1(n564), .A2(f[0]), .ZN(n578) );
  NAND2_X1 U487 ( .A1(n390), .A2(n389), .ZN(n590) );
  OAI21_X1 U488 ( .B1(n589), .B2(n593), .A(n590), .ZN(n586) );
  AOI21_X1 U489 ( .B1(n584), .B2(n586), .A(n582), .ZN(n606) );
  XNOR2_X1 U490 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U491 ( .A(n396), .B(n395), .ZN(n406) );
  INV_X1 U492 ( .A(n402), .ZN(n397) );
  NAND2_X1 U493 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U494 ( .A1(n406), .A2(n405), .ZN(n603) );
  OAI21_X1 U495 ( .B1(n606), .B2(n602), .A(n603), .ZN(n599) );
  OR2_X1 U496 ( .A1(n408), .A2(n407), .ZN(n597) );
  NAND2_X1 U497 ( .A1(n599), .A2(n597), .ZN(n609) );
  OAI22_X1 U498 ( .A1(n412), .A2(n411), .B1(n410), .B2(n409), .ZN(n445) );
  OAI22_X1 U499 ( .A1(n95), .A2(n415), .B1(n414), .B2(n413), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n649), .B(a_in[6]), .ZN(n436) );
  OAI22_X1 U501 ( .A1(n437), .A2(n418), .B1(n436), .B2(n689), .ZN(n439) );
  INV_X1 U502 ( .A(n170), .ZN(n419) );
  AND2_X1 U503 ( .A1(a_in[0]), .A2(n419), .ZN(n438) );
  FA_X1 U504 ( .A(n422), .B(n421), .CI(n420), .CO(n449), .S(n427) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n423) );
  XNOR2_X1 U506 ( .A(n448), .B(n423), .ZN(n433) );
  NAND2_X1 U507 ( .A1(n433), .A2(n432), .ZN(n613) );
  NAND3_X1 U508 ( .A1(n596), .A2(n609), .A3(n613), .ZN(n453) );
  HA_X1 U509 ( .A(n434), .B(f[7]), .CO(n461), .S(n468) );
  OAI22_X1 U510 ( .A1(n437), .A2(n436), .B1(n435), .B2(n689), .ZN(n467) );
  FA_X1 U511 ( .A(n439), .B(f[6]), .CI(n438), .CO(n466), .S(n450) );
  FA_X1 U512 ( .A(n440), .B(n441), .CI(n442), .CO(n462), .S(n484) );
  FA_X1 U513 ( .A(n445), .B(n444), .CI(n443), .CO(n483), .S(n448) );
  XNOR2_X1 U514 ( .A(n484), .B(n483), .ZN(n446) );
  XNOR2_X1 U515 ( .A(n482), .B(n446), .ZN(n455) );
  OR2_X1 U516 ( .A1(n449), .A2(n450), .ZN(n447) );
  NAND2_X1 U517 ( .A1(n450), .A2(n449), .ZN(n451) );
  OR2_X1 U518 ( .A1(n455), .A2(n454), .ZN(n617) );
  NAND3_X1 U519 ( .A1(n453), .A2(n615), .A3(n617), .ZN(n456) );
  NAND2_X1 U520 ( .A1(n455), .A2(n454), .ZN(n616) );
  NAND2_X1 U521 ( .A1(n456), .A2(n616), .ZN(n623) );
  XNOR2_X1 U522 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U523 ( .A(n460), .B(n459), .ZN(n490) );
  XNOR2_X1 U524 ( .A(n462), .B(n461), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(n464), .ZN(n478) );
  FA_X1 U526 ( .A(n466), .B(n467), .CI(n468), .CO(n476), .S(n482) );
  FA_X1 U527 ( .A(n471), .B(n470), .CI(n469), .CO(n306), .S(n475) );
  OR2_X1 U528 ( .A1(n476), .A2(n475), .ZN(n472) );
  NAND2_X1 U529 ( .A1(n478), .A2(n472), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n473), .ZN(n489) );
  XNOR2_X1 U532 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n478), .B(n477), .ZN(n488) );
  NOR2_X1 U534 ( .A1(n103), .A2(n628), .ZN(n536) );
  NAND2_X1 U535 ( .A1(n488), .A2(n487), .ZN(n627) );
  NAND2_X1 U536 ( .A1(n490), .A2(n489), .ZN(n630) );
  OAI21_X1 U537 ( .B1(n102), .B2(n627), .A(n630), .ZN(n535) );
  NOR2_X1 U538 ( .A1(n492), .A2(n491), .ZN(n518) );
  NOR2_X1 U539 ( .A1(n493), .A2(n494), .ZN(n520) );
  NOR2_X1 U540 ( .A1(n518), .A2(n520), .ZN(n496) );
  NAND2_X1 U541 ( .A1(n495), .A2(n496), .ZN(n538) );
  NOR2_X1 U542 ( .A1(n539), .A2(n538), .ZN(n497) );
  NAND2_X1 U543 ( .A1(n497), .A2(n126), .ZN(n502) );
  NOR2_X1 U544 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND3_X1 U545 ( .A1(n501), .A2(n502), .A3(n500), .ZN(n507) );
  INV_X1 U546 ( .A(n502), .ZN(n504) );
  NAND2_X1 U547 ( .A1(n504), .A2(n498), .ZN(n505) );
  NAND4_X1 U548 ( .A1(n508), .A2(n507), .A3(n506), .A4(n505), .ZN(n509) );
  NOR2_X2 U549 ( .A1(enable_f), .A2(reset), .ZN(n662) );
  NAND2_X1 U550 ( .A1(n509), .A2(n131), .ZN(n48) );
  INV_X1 U551 ( .A(n657), .ZN(n640) );
  OR2_X1 U552 ( .A1(n92), .A2(n518), .ZN(n656) );
  INV_X1 U553 ( .A(n656), .ZN(n512) );
  INV_X1 U554 ( .A(n510), .ZN(n654) );
  INV_X1 U555 ( .A(n654), .ZN(n511) );
  AOI21_X1 U556 ( .B1(n640), .B2(n512), .A(n511), .ZN(n515) );
  INV_X1 U557 ( .A(n110), .ZN(n513) );
  NAND2_X1 U558 ( .A1(n513), .A2(n101), .ZN(n514) );
  XNOR2_X1 U559 ( .A(n515), .B(n514), .ZN(n517) );
  NAND2_X1 U560 ( .A1(n662), .A2(f[12]), .ZN(n516) );
  OAI21_X1 U561 ( .B1(n517), .B2(n546), .A(n516), .ZN(n55) );
  INV_X1 U562 ( .A(n518), .ZN(n638) );
  INV_X1 U563 ( .A(n637), .ZN(n519) );
  AOI21_X1 U564 ( .B1(n640), .B2(n638), .A(n519), .ZN(n524) );
  INV_X1 U565 ( .A(n92), .ZN(n522) );
  NAND2_X1 U566 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U567 ( .A(n524), .B(n523), .ZN(n526) );
  NAND2_X1 U568 ( .A1(n662), .A2(f[11]), .ZN(n525) );
  OAI21_X1 U569 ( .B1(n526), .B2(n546), .A(n525), .ZN(n56) );
  OAI21_X1 U570 ( .B1(n657), .B2(n538), .A(n537), .ZN(n646) );
  OAI21_X1 U571 ( .B1(n554), .B2(n529), .A(n528), .ZN(n530) );
  AOI21_X1 U572 ( .B1(n646), .B2(n114), .A(n530), .ZN(n533) );
  XNOR2_X1 U573 ( .A(n533), .B(n117), .ZN(n534) );
  OAI21_X1 U574 ( .B1(n534), .B2(n546), .A(n127), .ZN(n49) );
  AOI21_X1 U575 ( .B1(n623), .B2(n536), .A(n535), .ZN(n539) );
  OAI21_X1 U576 ( .B1(n539), .B2(n538), .A(n537), .ZN(n557) );
  NOR2_X1 U577 ( .A1(n553), .A2(n540), .ZN(n542) );
  OAI21_X1 U578 ( .B1(n554), .B2(n540), .A(n558), .ZN(n541) );
  AOI21_X1 U579 ( .B1(n557), .B2(n542), .A(n541), .ZN(n545) );
  XNOR2_X1 U580 ( .A(n545), .B(n118), .ZN(n547) );
  INV_X1 U581 ( .A(n704), .ZN(n546) );
  OAI21_X1 U582 ( .B1(n547), .B2(n546), .A(n128), .ZN(n50) );
  AOI21_X1 U583 ( .B1(n557), .B2(n644), .A(n548), .ZN(n551) );
  XNOR2_X1 U584 ( .A(n551), .B(n119), .ZN(n552) );
  OAI21_X1 U585 ( .B1(n552), .B2(n546), .A(n129), .ZN(n52) );
  INV_X1 U586 ( .A(n553), .ZN(n556) );
  INV_X1 U587 ( .A(n554), .ZN(n555) );
  AOI21_X1 U588 ( .B1(n557), .B2(n556), .A(n555), .ZN(n560) );
  XNOR2_X1 U589 ( .A(n560), .B(n116), .ZN(n561) );
  OAI21_X1 U590 ( .B1(n561), .B2(n546), .A(n130), .ZN(n51) );
  INV_X1 U591 ( .A(n671), .ZN(n562) );
  OAI21_X1 U592 ( .B1(n691), .B2(n563), .A(n562), .ZN(n47) );
  OR2_X1 U593 ( .A1(n564), .A2(f[0]), .ZN(n565) );
  AND2_X1 U594 ( .A1(n565), .A2(n578), .ZN(n566) );
  AOI22_X1 U595 ( .A1(n566), .A2(n704), .B1(n662), .B2(f[0]), .ZN(n567) );
  INV_X1 U596 ( .A(n567), .ZN(n67) );
  NOR2_X2 U597 ( .A1(valid_in), .A2(reset), .ZN(n670) );
  AOI22_X1 U598 ( .A1(n671), .A2(b[0]), .B1(n670), .B2(b_in[0]), .ZN(n703) );
  AOI22_X1 U599 ( .A1(n671), .A2(a[9]), .B1(n670), .B2(a_in[9]), .ZN(n568) );
  INV_X1 U600 ( .A(n568), .ZN(n77) );
  AOI22_X1 U601 ( .A1(n671), .A2(a[8]), .B1(n670), .B2(a_in[8]), .ZN(n569) );
  INV_X1 U602 ( .A(n569), .ZN(n78) );
  AOI22_X1 U603 ( .A1(n671), .A2(a[7]), .B1(n670), .B2(a_in[7]), .ZN(n570) );
  INV_X1 U604 ( .A(n570), .ZN(n79) );
  AOI22_X1 U605 ( .A1(n671), .A2(a[6]), .B1(n670), .B2(a_in[6]), .ZN(n571) );
  INV_X1 U606 ( .A(n571), .ZN(n80) );
  AOI22_X1 U607 ( .A1(n671), .A2(a[5]), .B1(n670), .B2(a_in[5]), .ZN(n695) );
  AOI22_X1 U608 ( .A1(n671), .A2(a[0]), .B1(n670), .B2(a_in[0]), .ZN(n572) );
  INV_X1 U609 ( .A(n572), .ZN(n86) );
  AOI22_X1 U610 ( .A1(n671), .A2(a[4]), .B1(n670), .B2(a_in[4]), .ZN(n573) );
  INV_X1 U611 ( .A(n573), .ZN(n82) );
  AOI22_X1 U612 ( .A1(n671), .A2(a[3]), .B1(n670), .B2(a_in[3]), .ZN(n574) );
  INV_X1 U613 ( .A(n574), .ZN(n83) );
  AOI22_X1 U614 ( .A1(n671), .A2(a[2]), .B1(n670), .B2(a_in[2]), .ZN(n696) );
  AOI22_X1 U615 ( .A1(n671), .A2(a[1]), .B1(n670), .B2(a_in[1]), .ZN(n697) );
  AOI22_X1 U616 ( .A1(n671), .A2(b[8]), .B1(n670), .B2(b_in[8]), .ZN(n698) );
  AOI22_X1 U617 ( .A1(n671), .A2(b[2]), .B1(n670), .B2(b_in[2]), .ZN(n702) );
  AOI22_X1 U618 ( .A1(n671), .A2(b[4]), .B1(n670), .B2(b_in[4]), .ZN(n701) );
  NAND2_X1 U619 ( .A1(n124), .A2(n577), .ZN(n579) );
  XOR2_X1 U620 ( .A(n579), .B(n578), .Z(n580) );
  AOI22_X1 U621 ( .A1(n580), .A2(n704), .B1(n662), .B2(f[1]), .ZN(n581) );
  INV_X1 U622 ( .A(n581), .ZN(n66) );
  NAND2_X1 U623 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U624 ( .A(n100), .B(n585), .ZN(n587) );
  AOI22_X1 U625 ( .A1(n587), .A2(n704), .B1(n662), .B2(f[3]), .ZN(n588) );
  INV_X1 U626 ( .A(n588), .ZN(n64) );
  INV_X1 U627 ( .A(n589), .ZN(n591) );
  NAND2_X1 U628 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U629 ( .A(n593), .B(n592), .Z(n594) );
  AOI22_X1 U630 ( .A1(n594), .A2(n704), .B1(n662), .B2(f[2]), .ZN(n595) );
  INV_X1 U631 ( .A(n595), .ZN(n65) );
  NAND2_X1 U632 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U633 ( .A(n599), .B(n598), .ZN(n600) );
  AOI22_X1 U634 ( .A1(n600), .A2(n704), .B1(n662), .B2(f[5]), .ZN(n601) );
  INV_X1 U635 ( .A(n601), .ZN(n62) );
  INV_X1 U636 ( .A(n602), .ZN(n604) );
  NAND2_X1 U637 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U638 ( .A(n606), .B(n605), .Z(n607) );
  AOI22_X1 U639 ( .A1(n607), .A2(n704), .B1(n662), .B2(f[4]), .ZN(n608) );
  INV_X1 U640 ( .A(n608), .ZN(n63) );
  NAND2_X1 U641 ( .A1(n615), .A2(n613), .ZN(n610) );
  XNOR2_X1 U642 ( .A(n115), .B(n610), .ZN(n611) );
  AOI22_X1 U643 ( .A1(n611), .A2(n704), .B1(n662), .B2(f[6]), .ZN(n612) );
  INV_X1 U644 ( .A(n612), .ZN(n61) );
  INV_X1 U645 ( .A(n613), .ZN(n614) );
  AOI21_X1 U646 ( .B1(n115), .B2(n615), .A(n614), .ZN(n619) );
  NAND2_X1 U647 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U648 ( .A(n619), .B(n618), .Z(n620) );
  AOI22_X1 U649 ( .A1(n620), .A2(n704), .B1(n662), .B2(f[7]), .ZN(n621) );
  INV_X1 U650 ( .A(n621), .ZN(n60) );
  INV_X1 U651 ( .A(n628), .ZN(n622) );
  NAND2_X1 U652 ( .A1(n622), .A2(n627), .ZN(n624) );
  INV_X1 U653 ( .A(n99), .ZN(n629) );
  XOR2_X1 U654 ( .A(n624), .B(n629), .Z(n625) );
  AOI22_X1 U655 ( .A1(n625), .A2(n704), .B1(n662), .B2(f[8]), .ZN(n626) );
  INV_X1 U656 ( .A(n626), .ZN(n59) );
  OAI21_X1 U657 ( .B1(n629), .B2(n628), .A(n627), .ZN(n633) );
  INV_X1 U658 ( .A(n103), .ZN(n631) );
  NAND2_X1 U659 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U660 ( .A(n633), .B(n632), .ZN(n634) );
  NAND2_X1 U661 ( .A1(n634), .A2(n704), .ZN(n636) );
  NAND2_X1 U662 ( .A1(n662), .A2(f[9]), .ZN(n635) );
  NAND2_X1 U663 ( .A1(n636), .A2(n635), .ZN(n58) );
  NAND2_X1 U664 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U665 ( .A(n640), .B(n639), .ZN(n641) );
  AOI22_X1 U666 ( .A1(n641), .A2(n704), .B1(n662), .B2(f[10]), .ZN(n642) );
  INV_X1 U667 ( .A(n642), .ZN(n57) );
  NAND2_X1 U668 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U669 ( .A(n646), .B(n645), .ZN(n647) );
  AOI22_X1 U670 ( .A1(n647), .A2(n704), .B1(n662), .B2(f[14]), .ZN(n648) );
  INV_X1 U671 ( .A(n648), .ZN(n53) );
  AOI22_X1 U672 ( .A1(n671), .A2(b[6]), .B1(n670), .B2(b_in[6]), .ZN(n699) );
  AOI22_X1 U673 ( .A1(n671), .A2(b[1]), .B1(n670), .B2(n649), .ZN(n692) );
  AOI22_X1 U674 ( .A1(n671), .A2(b[9]), .B1(n670), .B2(n650), .ZN(n651) );
  INV_X1 U675 ( .A(n651), .ZN(n68) );
  AOI22_X1 U676 ( .A1(n671), .A2(b[3]), .B1(n670), .B2(n652), .ZN(n693) );
  AOI22_X1 U677 ( .A1(n671), .A2(b[7]), .B1(n670), .B2(n292), .ZN(n694) );
  OAI21_X1 U678 ( .B1(n654), .B2(n110), .A(n101), .ZN(n667) );
  NOR2_X1 U679 ( .A1(n125), .A2(n105), .ZN(n663) );
  OR2_X1 U680 ( .A1(n658), .A2(n109), .ZN(n661) );
  OR2_X1 U681 ( .A1(n663), .A2(n132), .ZN(n666) );
  AOI21_X1 U682 ( .B1(n123), .B2(n663), .A(n112), .ZN(n665) );
  NAND2_X1 U683 ( .A1(n667), .A2(n123), .ZN(n664) );
  OAI211_X1 U684 ( .C1(n667), .C2(n666), .A(n665), .B(n664), .ZN(n668) );
  AOI22_X1 U685 ( .A1(n671), .A2(b[5]), .B1(n670), .B2(n669), .ZN(n700) );
endmodule

